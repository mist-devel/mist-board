library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity rom16k is
    Port ( CLK : in  STD_LOGIC;
             A : in  STD_LOGIC_VECTOR (13 downto 0);
          DOUT : out STD_LOGIC_VECTOR (7 downto 0)
		   );
				
end rom16k;

architecture Behavioral of rom16k is

type
  -- 14K ROM 0000..37FF
  romarray is array(0 to 16383) of std_logic_vector(7 downto 0);

constant
  myROM : romarray := (

--x"f3",x"31",x"ff",x"7f",x"21",x"00",x"3c",x"11",x"01",x"3c",x"01",x"00",x"04",x"36",x"20",x"ed",
--x"b0",x"21",x"43",x"00",x"11",x"00",x"3e",x"cd",x"3b",x"00",x"21",x"55",x"00",x"11",x"80",x"3e",
--x"cd",x"3b",x"00",x"11",x"00",x"3c",x"21",x"01",x"38",x"4e",x"06",x"08",x"af",x"cb",x"01",x"ce",
--x"00",x"12",x"1c",x"10",x"f7",x"cb",x"05",x"30",x"f0",x"18",x"e8",x"7e",x"b7",x"c8",x"23",x"12",
--x"13",x"18",x"f8",x"48",x"54",x"31",x"30",x"38",x"30",x"5a",x"20",x"74",x"65",x"73",x"74",x"20",
--x"63",x"6f",x"64",x"65",x"00",x"41",x"6e",x"6f",x"74",x"68",x"65",x"72",x"20",x"74",x"65",x"73",
--x"74",x"20",x"74",x"65",x"78",x"74",x"2e",x"20",x"48",x"65",x"6c",x"6c",x"6f",x"20",x"77",x"6f",
--x"72",x"6c",x"64",x"21",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

--x"f3",x"31",x"ff",x"7f",x"21",x"00",x"3c",x"11",x"01",x"3c",x"01",x"00",x"04",x"36",x"20",x"ed",
--x"b0",x"af",x"21",x"00",x"3c",x"77",x"23",x"3c",x"20",x"fb",x"21",x"3a",x"00",x"11",x"00",x"3e",
--x"cd",x"32",x"00",x"21",x"4c",x"00",x"11",x"80",x"3e",x"cd",x"32",x"00",x"21",x"3f",x"3c",x"34",
--x"18",x"fd",x"7e",x"b7",x"c8",x"23",x"12",x"13",x"18",x"f8",x"48",x"54",x"31",x"30",x"38",x"30",
--x"5a",x"20",x"74",x"65",x"73",x"74",x"20",x"63",x"6f",x"64",x"65",x"00",x"41",x"6e",x"6f",x"74",
--x"68",x"65",x"72",x"20",x"74",x"65",x"73",x"74",x"20",x"74",x"65",x"78",x"74",x"2e",x"20",x"48",
--x"65",x"6c",x"6c",x"6f",x"20",x"77",x"6f",x"72",x"6c",x"64",x"21",x"00",x"00",x"00",x"00",x"00",

x"F3",x"AF",x"C3",x"74",x"06",x"C3",x"00",x"40",x"C3",x"00",x"40",x"E1",x"E9",x"C3",
x"9F",x"06",x"C3",x"03",x"40",x"C5",x"06",x"01",x"18",x"2E",x"C3",x"06",x"40",x"C5",
x"06",x"02",x"18",x"26",x"C3",x"09",x"40",x"C5",x"06",x"04",x"18",x"1E",x"C3",x"0C",
x"40",x"11",x"15",x"40",x"18",x"E3",x"C3",x"0F",x"40",x"11",x"1D",x"40",x"18",x"E3",
x"C3",x"12",x"40",x"11",x"25",x"40",x"18",x"DB",x"C3",x"D9",x"05",x"C9",x"00",x"00",
x"C3",x"C2",x"03",x"CD",x"2B",x"00",x"B7",x"C0",x"18",x"F9",x"0D",x"0D",x"1F",x"1F",
x"01",x"01",x"5B",x"1B",x"0A",x"1A",x"08",x"18",x"09",x"19",x"20",x"20",x"0B",x"78",
x"B1",x"20",x"FB",x"C9",x"31",x"00",x"06",x"3A",x"EC",x"37",x"3C",x"FE",x"02",x"D2",
x"00",x"00",x"C3",x"CC",x"06",x"11",x"80",x"40",x"21",x"F7",x"18",x"01",x"27",x"00",
x"ED",x"B0",x"21",x"E5",x"41",x"36",x"3A",x"23",x"70",x"23",x"36",x"2C",x"23",x"22",
x"A7",x"40",x"11",x"2D",x"01",x"06",x"1C",x"21",x"52",x"41",x"36",x"C3",x"23",x"73",
x"23",x"72",x"23",x"10",x"F7",x"06",x"15",x"36",x"C9",x"23",x"23",x"23",x"10",x"F9",
x"21",x"E8",x"42",x"70",x"31",x"F8",x"41",x"CD",x"8F",x"1B",x"CD",x"C9",x"01",x"21",
x"05",x"01",x"CD",x"A7",x"28",x"CD",x"B3",x"1B",x"38",x"F5",x"D7",x"B7",x"20",x"12",
x"21",x"4C",x"43",x"23",x"7C",x"B5",x"28",x"1B",x"7E",x"47",x"2F",x"77",x"BE",x"70",
x"28",x"F3",x"18",x"11",x"CD",x"5A",x"1E",x"B7",x"C2",x"97",x"19",x"EB",x"2B",x"3E",
x"8F",x"46",x"77",x"BE",x"70",x"20",x"CE",x"2B",x"11",x"14",x"44",x"DF",x"DA",x"7A",
x"19",x"11",x"CE",x"FF",x"22",x"B1",x"40",x"19",x"22",x"A0",x"40",x"CD",x"4D",x"1B",
x"21",x"11",x"01",x"CD",x"A7",x"28",x"C3",x"19",x"1A",x"52",x"45",x"41",x"44",x"59",
x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",
x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",
x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"00",x"1E",x"2C",x"C3",x"A2",x"19",x"D7",x"AF",
x"01",x"3E",x"80",x"01",x"3E",x"01",x"F5",x"CF",x"28",x"CD",x"1C",x"2B",x"FE",x"80",
x"D2",x"4A",x"1E",x"F5",x"CF",x"2C",x"CD",x"1C",x"2B",x"FE",x"30",x"D2",x"4A",x"1E",
x"16",x"FF",x"14",x"D6",x"03",x"30",x"FB",x"C6",x"03",x"4F",x"F1",x"87",x"5F",x"06",
x"02",x"7A",x"1F",x"57",x"7B",x"1F",x"5F",x"10",x"F8",x"79",x"8F",x"3C",x"47",x"AF",
x"37",x"8F",x"10",x"FD",x"4F",x"7A",x"F6",x"3C",x"57",x"1A",x"B7",x"FA",x"7C",x"01",
x"3E",x"80",x"47",x"F1",x"B7",x"78",x"28",x"10",x"12",x"FA",x"8F",x"01",x"79",x"2F",
x"4F",x"1A",x"A1",x"12",x"CF",x"29",x"C9",x"B1",x"18",x"F9",x"A1",x"C6",x"FF",x"9F",
x"E5",x"CD",x"8D",x"09",x"E1",x"18",x"EF",x"D7",x"E5",x"3A",x"99",x"40",x"B7",x"20",
x"06",x"CD",x"58",x"03",x"B7",x"28",x"11",x"F5",x"AF",x"32",x"99",x"40",x"3C",x"CD",
x"57",x"28",x"F1",x"2A",x"D4",x"40",x"77",x"C3",x"84",x"28",x"21",x"28",x"19",x"22",
x"21",x"41",x"3E",x"03",x"32",x"AF",x"40",x"E1",x"C9",x"3E",x"1C",x"CD",x"3A",x"03",
x"3E",x"1F",x"C3",x"3A",x"03",x"ED",x"5F",x"32",x"AB",x"40",x"C9",x"21",x"01",x"FC",
x"CD",x"21",x"02",x"06",x"0B",x"10",x"FE",x"21",x"02",x"FC",x"CD",x"21",x"02",x"06",
x"0B",x"10",x"FE",x"21",x"00",x"FC",x"CD",x"21",x"02",x"06",x"5C",x"10",x"FE",x"C9",
x"E5",x"21",x"00",x"FB",x"18",x"1B",x"7E",x"D6",x"23",x"3E",x"00",x"20",x"0D",x"CD",
x"01",x"2B",x"CF",x"2C",x"7B",x"A2",x"C6",x"02",x"D2",x"4A",x"1E",x"3D",x"D3",x"FE",
x"00",x"E5",x"21",x"04",x"FF",x"CD",x"21",x"02",x"E1",x"C9",x"21",x"00",x"FF",x"3A",
x"3D",x"40",x"A4",x"B5",x"D3",x"FF",x"32",x"3D",x"40",x"C9",x"3A",x"3F",x"3C",x"EE",
x"0A",x"32",x"3F",x"3C",x"C9",x"C5",x"E5",x"06",x"08",x"CD",x"41",x"02",x"10",x"FB",
x"E1",x"C1",x"C9",x"C5",x"F5",x"DB",x"FF",x"17",x"30",x"FB",x"06",x"41",x"10",x"FE",
x"CD",x"1E",x"02",x"06",x"76",x"10",x"FE",x"DB",x"FF",x"47",x"F1",x"CB",x"10",x"17",
x"F5",x"CD",x"1E",x"02",x"F1",x"C1",x"C9",x"CD",x"64",x"02",x"E5",x"C5",x"D5",x"F5",
x"0E",x"08",x"57",x"CD",x"D9",x"01",x"7A",x"07",x"57",x"30",x"0B",x"CD",x"D9",x"01",
x"0D",x"20",x"F2",x"F1",x"D1",x"C1",x"E1",x"C9",x"06",x"87",x"10",x"FE",x"18",x"F2",
x"CD",x"FE",x"01",x"06",x"FF",x"AF",x"CD",x"64",x"02",x"10",x"FB",x"3E",x"A5",x"18",
x"D1",x"CD",x"FE",x"01",x"E5",x"AF",x"CD",x"41",x"02",x"FE",x"A5",x"20",x"F9",x"3E",
x"2A",x"32",x"3E",x"3C",x"32",x"3F",x"3C",x"E1",x"C9",x"CD",x"14",x"03",x"22",x"DF",
x"40",x"CD",x"F8",x"01",x"CD",x"E2",x"41",x"31",x"88",x"42",x"CD",x"FE",x"20",x"3E",
x"2A",x"CD",x"2A",x"03",x"CD",x"B3",x"1B",x"DA",x"CC",x"06",x"D7",x"CA",x"97",x"19",
x"FE",x"2F",x"28",x"4F",x"CD",x"93",x"02",x"CD",x"35",x"02",x"FE",x"55",x"20",x"F9",
x"06",x"06",x"7E",x"B7",x"28",x"09",x"CD",x"35",x"02",x"BE",x"20",x"ED",x"23",x"10",
x"F3",x"CD",x"2C",x"02",x"CD",x"35",x"02",x"FE",x"78",x"28",x"B8",x"FE",x"3C",x"20",
x"F5",x"CD",x"35",x"02",x"47",x"CD",x"14",x"03",x"85",x"4F",x"CD",x"35",x"02",x"77",
x"23",x"81",x"4F",x"10",x"F7",x"CD",x"35",x"02",x"B9",x"28",x"DA",x"3E",x"43",x"32",
x"3E",x"3C",x"18",x"D6",x"CD",x"35",x"02",x"6F",x"CD",x"35",x"02",x"67",x"C9",x"EB",
x"2A",x"DF",x"40",x"EB",x"D7",x"C4",x"5A",x"1E",x"20",x"8A",x"EB",x"E9",x"C5",x"4F",
x"CD",x"C1",x"41",x"3A",x"9C",x"40",x"B7",x"79",x"C1",x"FA",x"64",x"02",x"20",x"62",
x"D5",x"CD",x"33",x"00",x"F5",x"CD",x"48",x"03",x"32",x"A6",x"40",x"F1",x"D1",x"C9",
x"3A",x"3D",x"40",x"E6",x"08",x"3A",x"20",x"40",x"28",x"03",x"0F",x"E6",x"1F",x"E6",
x"3F",x"C9",x"CD",x"C4",x"41",x"D5",x"CD",x"2B",x"00",x"D1",x"C9",x"AF",x"32",x"99",
x"40",x"32",x"A6",x"40",x"CD",x"AF",x"41",x"C5",x"2A",x"A7",x"40",x"06",x"F0",x"CD",
x"D9",x"05",x"F5",x"48",x"06",x"00",x"09",x"36",x"00",x"2A",x"A7",x"40",x"F1",x"C1",
x"2B",x"D8",x"AF",x"C9",x"CD",x"58",x"03",x"B7",x"C0",x"18",x"F9",x"AF",x"32",x"9C",
x"40",x"3A",x"9B",x"40",x"B7",x"C8",x"3E",x"0D",x"D5",x"CD",x"9C",x"03",x"D1",x"C9",
x"F5",x"D5",x"C5",x"4F",x"1E",x"00",x"FE",x"0C",x"28",x"10",x"FE",x"0A",x"20",x"03",
x"3E",x"0D",x"4F",x"FE",x"0D",x"28",x"05",x"3A",x"9B",x"40",x"3C",x"5F",x"7B",x"32",
x"9B",x"40",x"79",x"CD",x"3B",x"00",x"C1",x"D1",x"F1",x"C9",x"E5",x"DD",x"E5",x"D5",
x"DD",x"E1",x"D5",x"21",x"DD",x"03",x"E5",x"4F",x"1A",x"A0",x"B8",x"C2",x"33",x"40",
x"FE",x"02",x"DD",x"6E",x"01",x"DD",x"66",x"02",x"E9",x"D1",x"DD",x"E1",x"E1",x"C1",
x"C9",x"21",x"36",x"40",x"01",x"01",x"38",x"16",x"00",x"0A",x"5F",x"AE",x"73",x"A3",
x"20",x"08",x"14",x"2C",x"CB",x"01",x"F2",x"EB",x"03",x"C9",x"5F",x"7A",x"07",x"07",
x"07",x"57",x"0E",x"01",x"79",x"A3",x"20",x"05",x"14",x"CB",x"01",x"18",x"F7",x"3A",
x"80",x"38",x"47",x"7A",x"C6",x"40",x"FE",x"60",x"30",x"13",x"CB",x"08",x"30",x"31",
x"C6",x"20",x"57",x"3A",x"40",x"38",x"E6",x"10",x"28",x"28",x"7A",x"D6",x"60",x"18",
x"22",x"D6",x"70",x"30",x"10",x"C6",x"40",x"FE",x"3C",x"38",x"02",x"EE",x"10",x"CB",
x"08",x"30",x"12",x"EE",x"10",x"18",x"0E",x"07",x"CB",x"08",x"30",x"01",x"3C",x"21",
x"50",x"00",x"4F",x"06",x"00",x"09",x"7E",x"57",x"01",x"AC",x"0D",x"CD",x"60",x"00",
x"7A",x"FE",x"01",x"C0",x"EF",x"C9",x"DD",x"6E",x"03",x"DD",x"66",x"04",x"38",x"3A",
x"DD",x"7E",x"05",x"B7",x"28",x"01",x"77",x"79",x"FE",x"20",x"DA",x"06",x"05",x"FE",
x"80",x"30",x"35",x"FE",x"40",x"38",x"08",x"D6",x"40",x"FE",x"20",x"38",x"02",x"D6",
x"20",x"CD",x"41",x"05",x"7C",x"E6",x"03",x"F6",x"3C",x"67",x"56",x"DD",x"7E",x"05",
x"B7",x"28",x"05",x"DD",x"72",x"05",x"36",x"5F",x"DD",x"75",x"03",x"DD",x"74",x"04",
x"79",x"C9",x"DD",x"7E",x"05",x"B7",x"C0",x"7E",x"C9",x"7D",x"E6",x"C0",x"6F",x"C9",
x"FE",x"C0",x"38",x"D3",x"D6",x"C0",x"28",x"D2",x"47",x"3E",x"20",x"CD",x"41",x"05",
x"10",x"F9",x"18",x"C8",x"7E",x"DD",x"77",x"05",x"C9",x"AF",x"18",x"F9",x"21",x"00",
x"3C",x"3A",x"3D",x"40",x"E6",x"F7",x"32",x"3D",x"40",x"D3",x"FF",x"C9",x"2B",x"3A",
x"3D",x"40",x"E6",x"08",x"28",x"01",x"2B",x"36",x"20",x"C9",x"3A",x"3D",x"40",x"E6",
x"08",x"C4",x"E2",x"04",x"7D",x"E6",x"3F",x"2B",x"C0",x"11",x"40",x"00",x"19",x"C9",
x"23",x"7D",x"E6",x"3F",x"C0",x"11",x"C0",x"FF",x"19",x"C9",x"3A",x"3D",x"40",x"F6",
x"08",x"32",x"3D",x"40",x"D3",x"FF",x"23",x"7D",x"E6",x"FE",x"6F",x"C9",x"11",x"80",
x"04",x"D5",x"FE",x"08",x"28",x"C0",x"FE",x"0A",x"D8",x"FE",x"0E",x"38",x"4F",x"28",
x"A1",x"FE",x"0F",x"28",x"A2",x"FE",x"17",x"28",x"D7",x"FE",x"18",x"28",x"B7",x"FE",
x"19",x"28",x"C5",x"FE",x"1A",x"28",x"BC",x"FE",x"1B",x"28",x"C2",x"FE",x"1C",x"28",
x"8D",x"FE",x"1D",x"CA",x"A1",x"04",x"FE",x"1E",x"28",x"37",x"FE",x"1F",x"28",x"3C",
x"C9",x"77",x"23",x"3A",x"3D",x"40",x"E6",x"08",x"28",x"01",x"23",x"7C",x"FE",x"40",
x"C0",x"11",x"C0",x"FF",x"19",x"E5",x"11",x"00",x"3C",x"21",x"40",x"3C",x"C5",x"01",
x"C0",x"03",x"ED",x"B0",x"C1",x"EB",x"18",x"19",x"7D",x"E6",x"C0",x"6F",x"E5",x"11",
x"40",x"00",x"19",x"7C",x"FE",x"40",x"28",x"E2",x"D1",x"E5",x"54",x"7D",x"F6",x"3F",
x"5F",x"13",x"18",x"04",x"E5",x"11",x"00",x"40",x"36",x"20",x"23",x"7C",x"BA",x"20",
x"F9",x"7D",x"BB",x"20",x"F5",x"E1",x"C9",x"79",x"B7",x"28",x"40",x"FE",x"0B",x"28",
x"0A",x"FE",x"0C",x"20",x"1B",x"AF",x"DD",x"B6",x"03",x"28",x"15",x"DD",x"7E",x"03",
x"DD",x"96",x"04",x"47",x"CD",x"D1",x"05",x"20",x"FB",x"3E",x"0A",x"00",x"D3",x"FD",
x"10",x"F4",x"18",x"18",x"F5",x"CD",x"D1",x"05",x"20",x"FB",x"F1",x"00",x"D3",x"FD",
x"FE",x"0D",x"C0",x"DD",x"34",x"04",x"DD",x"7E",x"04",x"DD",x"BE",x"03",x"79",x"C0",
x"DD",x"36",x"04",x"00",x"C9",x"00",x"DB",x"FD",x"E6",x"F0",x"FE",x"30",x"C9",x"E5",
x"3E",x"0E",x"CD",x"33",x"00",x"48",x"CD",x"49",x"00",x"FE",x"20",x"30",x"25",x"FE",
x"0D",x"CA",x"62",x"06",x"FE",x"1F",x"28",x"29",x"FE",x"01",x"28",x"6D",x"11",x"E0",
x"05",x"D5",x"FE",x"08",x"28",x"34",x"FE",x"18",x"28",x"2B",x"FE",x"09",x"28",x"42",
x"FE",x"19",x"28",x"39",x"FE",x"0A",x"C0",x"D1",x"77",x"78",x"B7",x"28",x"CF",x"7E",
x"23",x"CD",x"33",x"00",x"05",x"18",x"C7",x"CD",x"C9",x"01",x"41",x"E1",x"E5",x"C3",
x"E0",x"05",x"CD",x"30",x"06",x"2B",x"7E",x"23",x"FE",x"0A",x"C8",x"78",x"B9",x"20",
x"F3",x"C9",x"78",x"B9",x"C8",x"2B",x"7E",x"FE",x"0A",x"23",x"C8",x"2B",x"3E",x"08",
x"CD",x"33",x"00",x"04",x"C9",x"3E",x"17",x"C3",x"33",x"00",x"CD",x"48",x"03",x"E6",
x"07",x"2F",x"3C",x"C6",x"08",x"5F",x"78",x"B7",x"C8",x"3E",x"20",x"77",x"23",x"D5",
x"CD",x"33",x"00",x"D1",x"05",x"1D",x"C8",x"18",x"EF",x"37",x"F5",x"3E",x"0D",x"77",
x"CD",x"33",x"00",x"3E",x"0F",x"CD",x"33",x"00",x"79",x"90",x"47",x"F1",x"E1",x"C9",
x"D3",x"FF",x"21",x"D2",x"06",x"11",x"00",x"40",x"01",x"36",x"00",x"ED",x"B0",x"3D",
x"3D",x"20",x"F1",x"06",x"27",x"12",x"13",x"10",x"FC",x"3A",x"40",x"38",x"E6",x"04",
x"C2",x"75",x"00",x"31",x"7D",x"40",x"3A",x"EC",x"37",x"3C",x"FE",x"02",x"DA",x"75",
x"00",x"3E",x"01",x"32",x"E1",x"37",x"21",x"EC",x"37",x"11",x"EF",x"37",x"36",x"03",
x"01",x"00",x"00",x"CD",x"60",x"00",x"CB",x"46",x"20",x"FC",x"AF",x"32",x"EE",x"37",
x"01",x"00",x"42",x"3E",x"8C",x"77",x"CB",x"4E",x"28",x"FC",x"1A",x"02",x"0C",x"20",
x"F7",x"C3",x"00",x"42",x"01",x"18",x"1A",x"C3",x"AE",x"19",x"C3",x"96",x"1C",x"C3",
x"78",x"1D",x"C3",x"90",x"1C",x"C3",x"D9",x"25",x"C9",x"00",x"00",x"C9",x"00",x"00",
x"FB",x"C9",x"00",x"01",x"E3",x"03",x"00",x"00",x"00",x"4B",x"49",x"07",x"58",x"04",
x"00",x"3C",x"00",x"44",x"4F",x"06",x"8D",x"05",x"43",x"00",x"00",x"50",x"52",x"C3",
x"00",x"50",x"C7",x"00",x"00",x"3E",x"00",x"C9",x"21",x"80",x"13",x"CD",x"C2",x"09",
x"18",x"06",x"CD",x"C2",x"09",x"CD",x"82",x"09",x"78",x"B7",x"C8",x"3A",x"24",x"41",
x"B7",x"CA",x"B4",x"09",x"90",x"30",x"0C",x"2F",x"3C",x"EB",x"CD",x"A4",x"09",x"EB",
x"CD",x"B4",x"09",x"C1",x"D1",x"FE",x"19",x"D0",x"F5",x"CD",x"DF",x"09",x"67",x"F1",
x"CD",x"D7",x"07",x"B4",x"21",x"21",x"41",x"F2",x"54",x"07",x"CD",x"B7",x"07",x"D2",
x"96",x"07",x"23",x"34",x"CA",x"B2",x"07",x"2E",x"01",x"CD",x"EB",x"07",x"18",x"42",
x"AF",x"90",x"47",x"7E",x"9B",x"5F",x"23",x"7E",x"9A",x"57",x"23",x"7E",x"99",x"4F",
x"DC",x"C3",x"07",x"68",x"63",x"AF",x"47",x"79",x"B7",x"20",x"18",x"4A",x"54",x"65",
x"6F",x"78",x"D6",x"08",x"FE",x"E0",x"20",x"F0",x"AF",x"32",x"24",x"41",x"C9",x"05",
x"29",x"7A",x"17",x"57",x"79",x"8F",x"4F",x"F2",x"7D",x"07",x"78",x"5C",x"45",x"B7",
x"28",x"08",x"21",x"24",x"41",x"86",x"77",x"30",x"E3",x"C8",x"78",x"21",x"24",x"41",
x"B7",x"FC",x"A8",x"07",x"46",x"23",x"7E",x"E6",x"80",x"A9",x"4F",x"C3",x"B4",x"09",
x"1C",x"C0",x"14",x"C0",x"0C",x"C0",x"0E",x"80",x"34",x"C0",x"1E",x"0A",x"C3",x"A2",
x"19",x"7E",x"83",x"5F",x"23",x"7E",x"8A",x"57",x"23",x"7E",x"89",x"4F",x"C9",x"21",
x"25",x"41",x"7E",x"2F",x"77",x"AF",x"6F",x"90",x"47",x"7D",x"9B",x"5F",x"7D",x"9A",
x"57",x"7D",x"99",x"4F",x"C9",x"06",x"00",x"D6",x"08",x"38",x"07",x"43",x"5A",x"51",
x"0E",x"00",x"18",x"F5",x"C6",x"09",x"6F",x"AF",x"2D",x"C8",x"79",x"1F",x"4F",x"7A",
x"1F",x"57",x"7B",x"1F",x"5F",x"78",x"1F",x"47",x"18",x"EF",x"00",x"00",x"00",x"81",
x"03",x"AA",x"56",x"19",x"80",x"F1",x"22",x"76",x"80",x"45",x"AA",x"38",x"82",x"CD",
x"55",x"09",x"B7",x"EA",x"4A",x"1E",x"21",x"24",x"41",x"7E",x"01",x"35",x"80",x"11",
x"F3",x"04",x"90",x"F5",x"70",x"D5",x"C5",x"CD",x"16",x"07",x"C1",x"D1",x"04",x"CD",
x"A2",x"08",x"21",x"F8",x"07",x"CD",x"10",x"07",x"21",x"FC",x"07",x"CD",x"9A",x"14",
x"01",x"80",x"80",x"11",x"00",x"00",x"CD",x"16",x"07",x"F1",x"CD",x"89",x"0F",x"01",
x"31",x"80",x"11",x"18",x"72",x"CD",x"55",x"09",x"C8",x"2E",x"00",x"CD",x"14",x"09",
x"79",x"32",x"4F",x"41",x"EB",x"22",x"50",x"41",x"01",x"00",x"00",x"50",x"58",x"21",
x"65",x"07",x"E5",x"21",x"69",x"08",x"E5",x"E5",x"21",x"21",x"41",x"7E",x"23",x"B7",
x"28",x"24",x"E5",x"2E",x"08",x"1F",x"67",x"79",x"30",x"0B",x"E5",x"2A",x"50",x"41",
x"19",x"EB",x"E1",x"3A",x"4F",x"41",x"89",x"1F",x"4F",x"7A",x"1F",x"57",x"7B",x"1F",
x"5F",x"78",x"1F",x"47",x"2D",x"7C",x"20",x"E1",x"E1",x"C9",x"43",x"5A",x"51",x"4F",
x"C9",x"CD",x"A4",x"09",x"21",x"D8",x"0D",x"CD",x"B1",x"09",x"C1",x"D1",x"CD",x"55",
x"09",x"CA",x"9A",x"19",x"2E",x"FF",x"CD",x"14",x"09",x"34",x"34",x"2B",x"7E",x"32",
x"89",x"40",x"2B",x"7E",x"32",x"85",x"40",x"2B",x"7E",x"32",x"81",x"40",x"41",x"EB",
x"AF",x"4F",x"57",x"5F",x"32",x"8C",x"40",x"E5",x"C5",x"7D",x"CD",x"80",x"40",x"DE",
x"00",x"3F",x"30",x"07",x"32",x"8C",x"40",x"F1",x"F1",x"37",x"D2",x"C1",x"E1",x"79",
x"3C",x"3D",x"1F",x"FA",x"97",x"07",x"17",x"7B",x"17",x"5F",x"7A",x"17",x"57",x"79",
x"17",x"4F",x"29",x"78",x"17",x"47",x"3A",x"8C",x"40",x"17",x"32",x"8C",x"40",x"79",
x"B2",x"B3",x"20",x"CB",x"E5",x"21",x"24",x"41",x"35",x"E1",x"20",x"C3",x"C3",x"B2",
x"07",x"3E",x"FF",x"2E",x"AF",x"21",x"2D",x"41",x"4E",x"23",x"AE",x"47",x"2E",x"00",
x"78",x"B7",x"28",x"1F",x"7D",x"21",x"24",x"41",x"AE",x"80",x"47",x"1F",x"A8",x"78",
x"F2",x"36",x"09",x"C6",x"80",x"77",x"CA",x"90",x"08",x"CD",x"DF",x"09",x"77",x"2B",
x"C9",x"CD",x"55",x"09",x"2F",x"E1",x"B7",x"E1",x"F2",x"78",x"07",x"C3",x"B2",x"07",
x"CD",x"BF",x"09",x"78",x"B7",x"C8",x"C6",x"02",x"DA",x"B2",x"07",x"47",x"CD",x"16",
x"07",x"21",x"24",x"41",x"34",x"C0",x"C3",x"B2",x"07",x"3A",x"24",x"41",x"B7",x"C8",
x"3A",x"23",x"41",x"FE",x"2F",x"17",x"9F",x"C0",x"3C",x"C9",x"06",x"88",x"11",x"00",
x"00",x"21",x"24",x"41",x"4F",x"70",x"06",x"00",x"23",x"36",x"80",x"17",x"C3",x"62",
x"07",x"CD",x"94",x"09",x"F0",x"E7",x"FA",x"5B",x"0C",x"CA",x"F6",x"0A",x"21",x"23",
x"41",x"7E",x"EE",x"80",x"77",x"C9",x"CD",x"94",x"09",x"6F",x"17",x"9F",x"67",x"C3",
x"9A",x"0A",x"E7",x"CA",x"F6",x"0A",x"F2",x"55",x"09",x"2A",x"21",x"41",x"7C",x"B5",
x"C8",x"7C",x"18",x"BB",x"EB",x"2A",x"21",x"41",x"E3",x"E5",x"2A",x"23",x"41",x"E3",
x"E5",x"EB",x"C9",x"CD",x"C2",x"09",x"EB",x"22",x"21",x"41",x"60",x"69",x"22",x"23",
x"41",x"EB",x"C9",x"21",x"21",x"41",x"5E",x"23",x"56",x"23",x"4E",x"23",x"46",x"23",
x"C9",x"11",x"21",x"41",x"06",x"04",x"18",x"05",x"EB",x"3A",x"AF",x"40",x"47",x"1A",
x"77",x"13",x"23",x"05",x"20",x"F9",x"C9",x"21",x"23",x"41",x"7E",x"07",x"37",x"1F",
x"77",x"3F",x"1F",x"23",x"23",x"77",x"79",x"07",x"37",x"1F",x"4F",x"1F",x"AE",x"C9",
x"21",x"27",x"41",x"11",x"D2",x"09",x"18",x"06",x"21",x"27",x"41",x"11",x"D3",x"09",
x"D5",x"11",x"21",x"41",x"E7",x"D8",x"11",x"1D",x"41",x"C9",x"78",x"B7",x"CA",x"55",
x"09",x"21",x"5E",x"09",x"E5",x"CD",x"55",x"09",x"79",x"C8",x"21",x"23",x"41",x"AE",
x"79",x"F8",x"CD",x"26",x"0A",x"1F",x"A9",x"C9",x"23",x"78",x"BE",x"C0",x"2B",x"79",
x"BE",x"C0",x"2B",x"7A",x"BE",x"C0",x"2B",x"7B",x"96",x"C0",x"E1",x"E1",x"C9",x"7A",
x"AC",x"7C",x"FA",x"5F",x"09",x"BA",x"C2",x"60",x"09",x"7D",x"93",x"C2",x"60",x"09",
x"C9",x"21",x"27",x"41",x"CD",x"D3",x"09",x"11",x"2E",x"41",x"1A",x"B7",x"CA",x"55",
x"09",x"21",x"5E",x"09",x"E5",x"CD",x"55",x"09",x"1B",x"1A",x"4F",x"C8",x"21",x"23",
x"41",x"AE",x"79",x"F8",x"13",x"23",x"06",x"08",x"1A",x"96",x"C2",x"23",x"0A",x"1B",
x"2B",x"05",x"20",x"F6",x"C1",x"C9",x"CD",x"4F",x"0A",x"C2",x"5E",x"09",x"C9",x"E7",
x"2A",x"21",x"41",x"F8",x"CA",x"F6",x"0A",x"D4",x"B9",x"0A",x"21",x"B2",x"07",x"E5",
x"3A",x"24",x"41",x"FE",x"90",x"30",x"0E",x"CD",x"FB",x"0A",x"EB",x"D1",x"22",x"21",
x"41",x"3E",x"02",x"32",x"AF",x"40",x"C9",x"01",x"80",x"90",x"11",x"00",x"00",x"CD",
x"0C",x"0A",x"C0",x"61",x"6A",x"18",x"E8",x"E7",x"E0",x"FA",x"CC",x"0A",x"CA",x"F6",
x"0A",x"CD",x"BF",x"09",x"CD",x"EF",x"0A",x"78",x"B7",x"C8",x"CD",x"DF",x"09",x"21",
x"20",x"41",x"46",x"C3",x"96",x"07",x"2A",x"21",x"41",x"CD",x"EF",x"0A",x"7C",x"55",
x"1E",x"00",x"06",x"90",x"C3",x"69",x"09",x"E7",x"D0",x"CA",x"F6",x"0A",x"FC",x"CC",
x"0A",x"21",x"00",x"00",x"22",x"1D",x"41",x"22",x"1F",x"41",x"3E",x"08",x"01",x"3E",
x"04",x"C3",x"9F",x"0A",x"E7",x"C8",x"1E",x"18",x"C3",x"A2",x"19",x"47",x"4F",x"57",
x"5F",x"B7",x"C8",x"E5",x"CD",x"BF",x"09",x"CD",x"DF",x"09",x"AE",x"67",x"FC",x"1F",
x"0B",x"3E",x"98",x"90",x"CD",x"D7",x"07",x"7C",x"17",x"DC",x"A8",x"07",x"06",x"00",
x"DC",x"C3",x"07",x"E1",x"C9",x"1B",x"7A",x"A3",x"3C",x"C0",x"0B",x"C9",x"E7",x"F8",
x"CD",x"55",x"09",x"F2",x"37",x"0B",x"CD",x"82",x"09",x"CD",x"37",x"0B",x"C3",x"7B",
x"09",x"E7",x"F8",x"30",x"1E",x"28",x"B9",x"CD",x"8E",x"0A",x"21",x"24",x"41",x"7E",
x"FE",x"98",x"3A",x"21",x"41",x"D0",x"7E",x"CD",x"FB",x"0A",x"36",x"98",x"7B",x"F5",
x"79",x"17",x"CD",x"62",x"07",x"F1",x"C9",x"21",x"24",x"41",x"7E",x"FE",x"90",x"DA",
x"7F",x"0A",x"20",x"14",x"4F",x"2B",x"7E",x"EE",x"80",x"06",x"06",x"2B",x"B6",x"05",
x"20",x"FB",x"B7",x"21",x"00",x"80",x"CA",x"9A",x"0A",x"79",x"FE",x"B8",x"D0",x"F5",
x"CD",x"BF",x"09",x"CD",x"DF",x"09",x"AE",x"2B",x"36",x"B8",x"F5",x"FC",x"A0",x"0B",
x"21",x"23",x"41",x"3E",x"B8",x"90",x"CD",x"69",x"0D",x"F1",x"FC",x"20",x"0D",x"AF",
x"32",x"1C",x"41",x"F1",x"D0",x"C3",x"D8",x"0C",x"21",x"1D",x"41",x"7E",x"35",x"B7",
x"23",x"28",x"FA",x"C9",x"E5",x"21",x"00",x"00",x"78",x"B1",x"28",x"12",x"3E",x"10",
x"29",x"DA",x"3D",x"27",x"EB",x"29",x"EB",x"30",x"04",x"09",x"DA",x"3D",x"27",x"3D",
x"20",x"F0",x"EB",x"E1",x"C9",x"7C",x"17",x"9F",x"47",x"CD",x"51",x"0C",x"79",x"98",
x"18",x"03",x"7C",x"17",x"9F",x"47",x"E5",x"7A",x"17",x"9F",x"19",x"88",x"0F",x"AC",
x"F2",x"99",x"0A",x"C5",x"EB",x"CD",x"CF",x"0A",x"F1",x"E1",x"CD",x"A4",x"09",x"EB",
x"CD",x"6B",x"0C",x"C3",x"8F",x"0F",x"7C",x"B5",x"CA",x"9A",x"0A",x"E5",x"D5",x"CD",
x"45",x"0C",x"C5",x"44",x"4D",x"21",x"00",x"00",x"3E",x"10",x"29",x"38",x"1F",x"EB",
x"29",x"EB",x"30",x"04",x"09",x"DA",x"26",x"0C",x"3D",x"20",x"F1",x"C1",x"D1",x"7C",
x"B7",x"FA",x"1F",x"0C",x"D1",x"78",x"C3",x"4D",x"0C",x"EE",x"80",x"B5",x"28",x"13",
x"EB",x"01",x"C1",x"E1",x"CD",x"CF",x"0A",x"E1",x"CD",x"A4",x"09",x"CD",x"CF",x"0A",
x"C1",x"D1",x"C3",x"47",x"08",x"78",x"B7",x"C1",x"FA",x"9A",x"0A",x"D5",x"CD",x"CF",
x"0A",x"D1",x"C3",x"82",x"09",x"7C",x"AA",x"47",x"CD",x"4C",x"0C",x"EB",x"7C",x"B7",
x"F2",x"9A",x"0A",x"AF",x"4F",x"95",x"6F",x"79",x"9C",x"67",x"C3",x"9A",x"0A",x"2A",
x"21",x"41",x"CD",x"51",x"0C",x"7C",x"EE",x"80",x"B5",x"C0",x"EB",x"CD",x"EF",x"0A",
x"AF",x"06",x"98",x"C3",x"69",x"09",x"21",x"2D",x"41",x"7E",x"EE",x"80",x"77",x"21",
x"2E",x"41",x"7E",x"B7",x"C8",x"47",x"2B",x"4E",x"11",x"24",x"41",x"1A",x"B7",x"CA",
x"F4",x"09",x"90",x"30",x"16",x"2F",x"3C",x"F5",x"0E",x"08",x"23",x"E5",x"1A",x"46",
x"77",x"78",x"12",x"1B",x"2B",x"0D",x"20",x"F6",x"E1",x"46",x"2B",x"4E",x"F1",x"FE",
x"39",x"D0",x"F5",x"CD",x"DF",x"09",x"23",x"36",x"00",x"47",x"F1",x"21",x"2D",x"41",
x"CD",x"69",x"0D",x"3A",x"26",x"41",x"32",x"1C",x"41",x"78",x"B7",x"F2",x"CF",x"0C",
x"CD",x"33",x"0D",x"D2",x"0E",x"0D",x"EB",x"34",x"CA",x"B2",x"07",x"CD",x"90",x"0D",
x"C3",x"0E",x"0D",x"CD",x"45",x"0D",x"21",x"25",x"41",x"DC",x"57",x"0D",x"AF",x"47",
x"3A",x"23",x"41",x"B7",x"20",x"1E",x"21",x"1C",x"41",x"0E",x"08",x"56",x"77",x"7A",
x"23",x"0D",x"20",x"F9",x"78",x"D6",x"08",x"FE",x"C0",x"20",x"E6",x"C3",x"78",x"07",
x"05",x"21",x"1C",x"41",x"CD",x"97",x"0D",x"B7",x"F2",x"F6",x"0C",x"78",x"B7",x"28",
x"09",x"21",x"24",x"41",x"86",x"77",x"D2",x"78",x"07",x"C8",x"3A",x"1C",x"41",x"B7",
x"FC",x"20",x"0D",x"21",x"25",x"41",x"7E",x"E6",x"80",x"2B",x"2B",x"AE",x"77",x"C9",
x"21",x"1D",x"41",x"06",x"07",x"34",x"C0",x"23",x"05",x"20",x"FA",x"34",x"CA",x"B2",
x"07",x"2B",x"36",x"80",x"C9",x"21",x"27",x"41",x"11",x"1D",x"41",x"0E",x"07",x"AF",
x"1A",x"8E",x"12",x"13",x"23",x"0D",x"20",x"F8",x"C9",x"21",x"27",x"41",x"11",x"1D",
x"41",x"0E",x"07",x"AF",x"1A",x"9E",x"12",x"13",x"23",x"0D",x"20",x"F8",x"C9",x"7E",
x"2F",x"77",x"21",x"1C",x"41",x"06",x"08",x"AF",x"4F",x"79",x"9E",x"77",x"23",x"05",
x"20",x"F9",x"C9",x"71",x"E5",x"D6",x"08",x"38",x"0E",x"E1",x"E5",x"11",x"00",x"08",
x"4E",x"73",x"59",x"2B",x"15",x"20",x"F9",x"18",x"EE",x"C6",x"09",x"57",x"AF",x"E1",
x"15",x"C8",x"E5",x"1E",x"08",x"7E",x"1F",x"77",x"2B",x"1D",x"20",x"F9",x"18",x"F0",
x"21",x"23",x"41",x"16",x"01",x"18",x"ED",x"0E",x"08",x"7E",x"17",x"77",x"23",x"0D",
x"20",x"F9",x"C9",x"CD",x"55",x"09",x"C8",x"CD",x"0A",x"09",x"CD",x"39",x"0E",x"71",
x"13",x"06",x"07",x"1A",x"13",x"B7",x"D5",x"28",x"17",x"0E",x"08",x"C5",x"1F",x"47",
x"DC",x"33",x"0D",x"CD",x"90",x"0D",x"78",x"C1",x"0D",x"20",x"F2",x"D1",x"05",x"20",
x"E6",x"C3",x"D8",x"0C",x"21",x"23",x"41",x"CD",x"70",x"0D",x"18",x"F1",x"00",x"00",
x"00",x"00",x"00",x"00",x"20",x"84",x"11",x"D4",x"0D",x"21",x"27",x"41",x"CD",x"D3",
x"09",x"3A",x"2E",x"41",x"B7",x"CA",x"9A",x"19",x"CD",x"07",x"09",x"34",x"34",x"CD",
x"39",x"0E",x"21",x"51",x"41",x"71",x"41",x"11",x"4A",x"41",x"21",x"27",x"41",x"CD",
x"4B",x"0D",x"1A",x"99",x"3F",x"38",x"0B",x"11",x"4A",x"41",x"21",x"27",x"41",x"CD",
x"39",x"0D",x"AF",x"DA",x"12",x"04",x"3A",x"23",x"41",x"3C",x"3D",x"1F",x"FA",x"11",
x"0D",x"17",x"21",x"1D",x"41",x"0E",x"07",x"CD",x"99",x"0D",x"21",x"4A",x"41",x"CD",
x"97",x"0D",x"78",x"B7",x"20",x"C9",x"21",x"24",x"41",x"35",x"20",x"C3",x"C3",x"B2",
x"07",x"79",x"32",x"2D",x"41",x"2B",x"11",x"50",x"41",x"01",x"00",x"07",x"7E",x"12",
x"71",x"1B",x"2B",x"05",x"20",x"F8",x"C9",x"CD",x"FC",x"09",x"EB",x"2B",x"7E",x"B7",
x"C8",x"C6",x"02",x"DA",x"B2",x"07",x"77",x"E5",x"CD",x"77",x"0C",x"E1",x"34",x"C0",
x"C3",x"B2",x"07",x"CD",x"78",x"07",x"CD",x"EC",x"0A",x"F6",x"AF",x"EB",x"01",x"FF",
x"00",x"60",x"68",x"CC",x"9A",x"0A",x"EB",x"7E",x"FE",x"2D",x"F5",x"CA",x"83",x"0E",
x"FE",x"2B",x"28",x"01",x"2B",x"D7",x"DA",x"29",x"0F",x"FE",x"2E",x"CA",x"E4",x"0E",
x"FE",x"45",x"28",x"14",x"FE",x"25",x"CA",x"EE",x"0E",x"FE",x"23",x"CA",x"F5",x"0E",
x"FE",x"21",x"CA",x"F6",x"0E",x"FE",x"44",x"20",x"24",x"B7",x"CD",x"FB",x"0E",x"E5",
x"21",x"BD",x"0E",x"E3",x"D7",x"15",x"FE",x"CE",x"C8",x"FE",x"2D",x"C8",x"14",x"FE",
x"CD",x"C8",x"FE",x"2B",x"C8",x"2B",x"F1",x"D7",x"DA",x"94",x"0F",x"14",x"20",x"03",
x"AF",x"93",x"5F",x"E5",x"7B",x"90",x"F4",x"0A",x"0F",x"FC",x"18",x"0F",x"20",x"F8",
x"E1",x"F1",x"E5",x"CC",x"7B",x"09",x"E1",x"E7",x"E8",x"E5",x"21",x"90",x"08",x"E5",
x"CD",x"A3",x"0A",x"C9",x"E7",x"0C",x"20",x"DF",x"DC",x"FB",x"0E",x"C3",x"83",x"0E",
x"E7",x"F2",x"97",x"19",x"23",x"18",x"D2",x"B7",x"CD",x"FB",x"0E",x"18",x"F7",x"E5",
x"D5",x"C5",x"F5",x"CC",x"B1",x"0A",x"F1",x"C4",x"DB",x"0A",x"C1",x"D1",x"E1",x"C9",
x"C8",x"F5",x"E7",x"F5",x"E4",x"3E",x"09",x"F1",x"EC",x"4D",x"0E",x"F1",x"3D",x"C9",
x"D5",x"E5",x"F5",x"E7",x"F5",x"E4",x"97",x"08",x"F1",x"EC",x"DC",x"0D",x"F1",x"E1",
x"D1",x"3C",x"C9",x"D5",x"78",x"89",x"47",x"C5",x"E5",x"7E",x"D6",x"30",x"F5",x"E7",
x"F2",x"5D",x"0F",x"2A",x"21",x"41",x"11",x"CD",x"0C",x"DF",x"30",x"19",x"54",x"5D",
x"29",x"29",x"19",x"29",x"F1",x"4F",x"09",x"7C",x"B7",x"FA",x"57",x"0F",x"22",x"21",
x"41",x"E1",x"C1",x"D1",x"C3",x"83",x"0E",x"79",x"F5",x"CD",x"CC",x"0A",x"37",x"30",
x"18",x"01",x"74",x"94",x"11",x"00",x"24",x"CD",x"0C",x"0A",x"F2",x"74",x"0F",x"CD",
x"3E",x"09",x"F1",x"CD",x"89",x"0F",x"18",x"DD",x"CD",x"E3",x"0A",x"CD",x"4D",x"0E",
x"CD",x"FC",x"09",x"F1",x"CD",x"64",x"09",x"CD",x"E3",x"0A",x"CD",x"77",x"0C",x"18",
x"C8",x"CD",x"A4",x"09",x"CD",x"64",x"09",x"C1",x"D1",x"C3",x"16",x"07",x"7B",x"FE",
x"0A",x"30",x"09",x"07",x"07",x"83",x"07",x"86",x"D6",x"30",x"5F",x"FA",x"1E",x"32",
x"C3",x"BD",x"0E",x"E5",x"21",x"24",x"19",x"CD",x"A7",x"28",x"E1",x"CD",x"9A",x"0A",
x"AF",x"CD",x"34",x"10",x"B6",x"CD",x"D9",x"0F",x"C3",x"A6",x"28",x"AF",x"CD",x"34",
x"10",x"E6",x"08",x"28",x"02",x"36",x"2B",x"EB",x"CD",x"94",x"09",x"EB",x"F2",x"D9",
x"0F",x"36",x"2D",x"C5",x"E5",x"CD",x"7B",x"09",x"E1",x"C1",x"B4",x"23",x"36",x"30",
x"3A",x"D8",x"40",x"57",x"17",x"3A",x"AF",x"40",x"DA",x"9A",x"10",x"CA",x"92",x"10",
x"FE",x"04",x"D2",x"3D",x"10",x"01",x"00",x"00",x"CD",x"2F",x"13",x"21",x"30",x"41",
x"46",x"0E",x"20",x"3A",x"D8",x"40",x"5F",x"E6",x"20",x"28",x"07",x"78",x"B9",x"0E",
x"2A",x"20",x"01",x"41",x"71",x"D7",x"28",x"14",x"FE",x"45",x"28",x"10",x"FE",x"44",
x"28",x"0C",x"FE",x"30",x"28",x"F0",x"FE",x"2C",x"28",x"EC",x"FE",x"2E",x"20",x"03",
x"2B",x"36",x"30",x"7B",x"E6",x"10",x"28",x"03",x"2B",x"36",x"24",x"7B",x"E6",x"04",
x"C0",x"2B",x"70",x"C9",x"32",x"D8",x"40",x"21",x"30",x"41",x"36",x"20",x"C9",x"FE",
x"05",x"E5",x"DE",x"00",x"17",x"57",x"14",x"CD",x"01",x"12",x"01",x"00",x"03",x"82",
x"FA",x"57",x"10",x"14",x"BA",x"30",x"04",x"3C",x"47",x"3E",x"02",x"D6",x"02",x"E1",
x"F5",x"CD",x"91",x"12",x"36",x"30",x"CC",x"C9",x"09",x"CD",x"A4",x"12",x"2B",x"7E",
x"FE",x"30",x"28",x"FA",x"FE",x"2E",x"C4",x"C9",x"09",x"F1",x"28",x"1F",x"F5",x"E7",
x"3E",x"22",x"8F",x"77",x"23",x"F1",x"36",x"2B",x"F2",x"85",x"10",x"36",x"2D",x"2F",
x"3C",x"06",x"2F",x"04",x"D6",x"0A",x"30",x"FB",x"C6",x"3A",x"23",x"70",x"23",x"77",
x"23",x"36",x"00",x"EB",x"21",x"30",x"41",x"C9",x"23",x"C5",x"FE",x"04",x"7A",x"D2",
x"09",x"11",x"1F",x"DA",x"A3",x"11",x"01",x"03",x"06",x"CD",x"89",x"12",x"D1",x"7A",
x"D6",x"05",x"F4",x"69",x"12",x"CD",x"2F",x"13",x"7B",x"B7",x"CC",x"2F",x"09",x"3D",
x"F4",x"69",x"12",x"E5",x"CD",x"F5",x"0F",x"E1",x"28",x"02",x"70",x"23",x"36",x"00",
x"21",x"2F",x"41",x"23",x"3A",x"F3",x"40",x"95",x"92",x"C8",x"7E",x"FE",x"20",x"28",
x"F4",x"FE",x"2A",x"28",x"F0",x"2B",x"E5",x"F5",x"01",x"DF",x"10",x"C5",x"D7",x"FE",
x"2D",x"C8",x"FE",x"2B",x"C8",x"FE",x"24",x"C8",x"C1",x"FE",x"30",x"20",x"0F",x"23",
x"D7",x"30",x"0B",x"2B",x"01",x"2B",x"77",x"F1",x"28",x"FB",x"C1",x"C3",x"CE",x"10",
x"F1",x"28",x"FD",x"E1",x"36",x"25",x"C9",x"E5",x"1F",x"DA",x"AA",x"11",x"28",x"14",
x"11",x"84",x"13",x"CD",x"49",x"0A",x"16",x"10",x"FA",x"32",x"11",x"E1",x"C1",x"CD",
x"BD",x"0F",x"2B",x"36",x"25",x"C9",x"01",x"0E",x"B6",x"11",x"CA",x"1B",x"CD",x"0C",
x"0A",x"F2",x"1B",x"11",x"16",x"06",x"CD",x"55",x"09",x"C4",x"01",x"12",x"E1",x"C1",
x"FA",x"57",x"11",x"C5",x"5F",x"78",x"92",x"93",x"F4",x"69",x"12",x"CD",x"7D",x"12",
x"CD",x"A4",x"12",x"B3",x"C4",x"77",x"12",x"B3",x"C4",x"91",x"12",x"D1",x"C3",x"B6",
x"10",x"5F",x"79",x"B7",x"C4",x"16",x"0F",x"83",x"FA",x"62",x"11",x"AF",x"C5",x"F5",
x"FC",x"18",x"0F",x"FA",x"64",x"11",x"C1",x"7B",x"90",x"C1",x"5F",x"82",x"78",x"FA",
x"7F",x"11",x"92",x"93",x"F4",x"69",x"12",x"C5",x"CD",x"7D",x"12",x"18",x"11",x"CD",
x"69",x"12",x"79",x"CD",x"94",x"12",x"4F",x"AF",x"92",x"93",x"CD",x"69",x"12",x"C5",
x"47",x"4F",x"CD",x"A4",x"12",x"C1",x"B1",x"20",x"03",x"2A",x"F3",x"40",x"83",x"3D",
x"F4",x"69",x"12",x"50",x"C3",x"BF",x"10",x"E5",x"D5",x"CD",x"CC",x"0A",x"D1",x"AF",
x"CA",x"B0",x"11",x"1E",x"10",x"01",x"1E",x"06",x"CD",x"55",x"09",x"37",x"C4",x"01",
x"12",x"E1",x"C1",x"F5",x"79",x"B7",x"F5",x"C4",x"16",x"0F",x"80",x"4F",x"7A",x"E6",
x"04",x"FE",x"01",x"9F",x"57",x"81",x"4F",x"93",x"F5",x"C5",x"FC",x"18",x"0F",x"FA",
x"D0",x"11",x"C1",x"F1",x"C5",x"F5",x"FA",x"DE",x"11",x"AF",x"2F",x"3C",x"80",x"3C",
x"82",x"47",x"0E",x"00",x"CD",x"A4",x"12",x"F1",x"F4",x"71",x"12",x"C1",x"F1",x"CC",
x"2F",x"09",x"F1",x"38",x"03",x"83",x"90",x"92",x"C5",x"CD",x"74",x"10",x"EB",x"D1",
x"C3",x"BF",x"10",x"D5",x"AF",x"F5",x"E7",x"E2",x"22",x"12",x"3A",x"24",x"41",x"FE",
x"91",x"D2",x"22",x"12",x"11",x"64",x"13",x"21",x"27",x"41",x"CD",x"D3",x"09",x"CD",
x"A1",x"0D",x"F1",x"D6",x"0A",x"F5",x"18",x"E6",x"CD",x"4F",x"12",x"E7",x"30",x"0B",
x"01",x"43",x"91",x"11",x"F9",x"4F",x"CD",x"0C",x"0A",x"18",x"06",x"11",x"6C",x"13",
x"CD",x"49",x"0A",x"F2",x"4B",x"12",x"F1",x"CD",x"0B",x"0F",x"F5",x"18",x"E2",x"F1",
x"CD",x"18",x"0F",x"F5",x"CD",x"4F",x"12",x"F1",x"B7",x"D1",x"C9",x"E7",x"EA",x"5E",
x"12",x"01",x"74",x"94",x"11",x"F8",x"23",x"CD",x"0C",x"0A",x"18",x"06",x"11",x"74",
x"13",x"CD",x"49",x"0A",x"E1",x"F2",x"43",x"12",x"E9",x"B7",x"C8",x"3D",x"36",x"30",
x"23",x"18",x"F9",x"20",x"04",x"C8",x"CD",x"91",x"12",x"36",x"30",x"23",x"3D",x"18",
x"F6",x"7B",x"82",x"3C",x"47",x"3C",x"D6",x"03",x"30",x"FC",x"C6",x"05",x"4F",x"3A",
x"D8",x"40",x"E6",x"40",x"C0",x"4F",x"C9",x"05",x"20",x"08",x"36",x"2E",x"22",x"F3",
x"40",x"23",x"48",x"C9",x"0D",x"C0",x"36",x"2C",x"23",x"0E",x"03",x"C9",x"D5",x"E7",
x"E2",x"EA",x"12",x"C5",x"E5",x"CD",x"FC",x"09",x"21",x"7C",x"13",x"CD",x"F7",x"09",
x"CD",x"77",x"0C",x"AF",x"CD",x"7B",x"0B",x"E1",x"C1",x"11",x"8C",x"13",x"3E",x"0A",
x"CD",x"91",x"12",x"C5",x"F5",x"E5",x"D5",x"06",x"2F",x"04",x"E1",x"E5",x"CD",x"48",
x"0D",x"30",x"F8",x"E1",x"CD",x"36",x"0D",x"EB",x"E1",x"70",x"23",x"F1",x"C1",x"3D",
x"20",x"E2",x"C5",x"E5",x"21",x"1D",x"41",x"CD",x"B1",x"09",x"18",x"0C",x"C5",x"E5",
x"CD",x"08",x"07",x"3C",x"CD",x"FB",x"0A",x"CD",x"B4",x"09",x"E1",x"C1",x"AF",x"11",
x"D2",x"13",x"3F",x"CD",x"91",x"12",x"C5",x"F5",x"E5",x"D5",x"CD",x"BF",x"09",x"E1",
x"06",x"2F",x"04",x"7B",x"96",x"5F",x"23",x"7A",x"9E",x"57",x"23",x"79",x"9E",x"4F",
x"2B",x"2B",x"30",x"F0",x"CD",x"B7",x"07",x"23",x"CD",x"B4",x"09",x"EB",x"E1",x"70",
x"23",x"F1",x"C1",x"38",x"D3",x"13",x"13",x"3E",x"04",x"18",x"06",x"D5",x"11",x"D8",
x"13",x"3E",x"05",x"CD",x"91",x"12",x"C5",x"F5",x"E5",x"EB",x"4E",x"23",x"46",x"C5",
x"23",x"E3",x"EB",x"2A",x"21",x"41",x"06",x"2F",x"04",x"7D",x"93",x"6F",x"7C",x"9A",
x"67",x"30",x"F7",x"19",x"22",x"21",x"41",x"D1",x"E1",x"70",x"23",x"F1",x"C1",x"3D",
x"20",x"D7",x"CD",x"91",x"12",x"77",x"D1",x"C9",x"00",x"00",x"00",x"00",x"F9",x"02",
x"15",x"A2",x"FD",x"FF",x"9F",x"31",x"A9",x"5F",x"63",x"B2",x"FE",x"FF",x"03",x"BF",
x"C9",x"1B",x"0E",x"B6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",
x"04",x"BF",x"C9",x"1B",x"0E",x"B6",x"00",x"80",x"C6",x"A4",x"7E",x"8D",x"03",x"00",
x"40",x"7A",x"10",x"F3",x"5A",x"00",x"00",x"A0",x"72",x"4E",x"18",x"09",x"00",x"00",
x"10",x"A5",x"D4",x"E8",x"00",x"00",x"00",x"E8",x"76",x"48",x"17",x"00",x"00",x"00",
x"E4",x"0B",x"54",x"02",x"00",x"00",x"00",x"CA",x"9A",x"3B",x"00",x"00",x"00",x"00",
x"E1",x"F5",x"05",x"00",x"00",x"00",x"80",x"96",x"98",x"00",x"00",x"00",x"00",x"40",
x"42",x"0F",x"00",x"00",x"00",x"00",x"A0",x"86",x"01",x"10",x"27",x"00",x"10",x"27",
x"E8",x"03",x"64",x"00",x"0A",x"00",x"01",x"00",x"21",x"82",x"09",x"E3",x"E9",x"CD",
x"A4",x"09",x"21",x"80",x"13",x"CD",x"B1",x"09",x"18",x"03",x"CD",x"B1",x"0A",x"C1",
x"D1",x"CD",x"55",x"09",x"78",x"28",x"3C",x"F2",x"04",x"14",x"B7",x"CA",x"9A",x"19",
x"B7",x"CA",x"79",x"07",x"D5",x"C5",x"79",x"F6",x"7F",x"CD",x"BF",x"09",x"F2",x"21",
x"14",x"D5",x"C5",x"CD",x"40",x"0B",x"C1",x"D1",x"F5",x"CD",x"0C",x"0A",x"E1",x"7C",
x"1F",x"E1",x"22",x"23",x"41",x"E1",x"22",x"21",x"41",x"DC",x"E2",x"13",x"CC",x"82",
x"09",x"D5",x"C5",x"CD",x"09",x"08",x"C1",x"D1",x"CD",x"47",x"08",x"CD",x"A4",x"09",
x"01",x"38",x"81",x"11",x"3B",x"AA",x"CD",x"47",x"08",x"3A",x"24",x"41",x"FE",x"88",
x"D2",x"31",x"09",x"CD",x"40",x"0B",x"C6",x"80",x"C6",x"02",x"DA",x"31",x"09",x"F5",
x"21",x"F8",x"07",x"CD",x"0B",x"07",x"CD",x"41",x"08",x"F1",x"C1",x"D1",x"F5",x"CD",
x"13",x"07",x"CD",x"82",x"09",x"21",x"79",x"14",x"CD",x"A9",x"14",x"11",x"00",x"00",
x"C1",x"4A",x"C3",x"47",x"08",x"08",x"40",x"2E",x"94",x"74",x"70",x"4F",x"2E",x"77",
x"6E",x"02",x"88",x"7A",x"E6",x"A0",x"2A",x"7C",x"50",x"AA",x"AA",x"7E",x"FF",x"FF",
x"7F",x"7F",x"00",x"00",x"80",x"81",x"00",x"00",x"00",x"81",x"CD",x"A4",x"09",x"11",
x"32",x"0C",x"D5",x"E5",x"CD",x"BF",x"09",x"CD",x"47",x"08",x"E1",x"CD",x"A4",x"09",
x"7E",x"23",x"CD",x"B1",x"09",x"06",x"F1",x"C1",x"D1",x"3D",x"C8",x"D5",x"C5",x"F5",
x"E5",x"CD",x"47",x"08",x"E1",x"CD",x"C2",x"09",x"E5",x"CD",x"16",x"07",x"E1",x"18",
x"E9",x"CD",x"7F",x"0A",x"7C",x"B7",x"FA",x"4A",x"1E",x"B5",x"CA",x"F0",x"14",x"E5",
x"CD",x"F0",x"14",x"CD",x"BF",x"09",x"EB",x"E3",x"C5",x"CD",x"CF",x"0A",x"C1",x"D1",
x"CD",x"47",x"08",x"21",x"F8",x"07",x"CD",x"0B",x"07",x"C3",x"40",x"0B",x"21",x"90",
x"40",x"E5",x"11",x"00",x"00",x"4B",x"26",x"03",x"2E",x"08",x"EB",x"29",x"EB",x"79",
x"17",x"4F",x"E3",x"7E",x"07",x"77",x"E3",x"D2",x"16",x"15",x"E5",x"2A",x"AA",x"40",
x"19",x"EB",x"3A",x"AC",x"40",x"89",x"4F",x"E1",x"2D",x"C2",x"FC",x"14",x"E3",x"23",
x"E3",x"25",x"C2",x"FA",x"14",x"E1",x"21",x"65",x"B0",x"19",x"22",x"AA",x"40",x"CD",
x"EF",x"0A",x"3E",x"05",x"89",x"32",x"AC",x"40",x"EB",x"06",x"80",x"21",x"25",x"41",
x"70",x"2B",x"70",x"4F",x"06",x"00",x"C3",x"65",x"07",x"21",x"8B",x"15",x"CD",x"0B",
x"07",x"CD",x"A4",x"09",x"01",x"49",x"83",x"11",x"DB",x"0F",x"CD",x"B4",x"09",x"C1",
x"D1",x"CD",x"A2",x"08",x"CD",x"A4",x"09",x"CD",x"40",x"0B",x"C1",x"D1",x"CD",x"13",
x"07",x"21",x"8F",x"15",x"CD",x"10",x"07",x"CD",x"55",x"09",x"37",x"F2",x"77",x"15",
x"CD",x"08",x"07",x"CD",x"55",x"09",x"B7",x"F5",x"F4",x"82",x"09",x"21",x"8F",x"15",
x"CD",x"0B",x"07",x"F1",x"D4",x"82",x"09",x"21",x"93",x"15",x"C3",x"9A",x"14",x"DB",
x"0F",x"49",x"81",x"00",x"00",x"00",x"7F",x"05",x"BA",x"D7",x"1E",x"86",x"64",x"26",
x"99",x"87",x"58",x"34",x"23",x"87",x"E0",x"5D",x"A5",x"86",x"DA",x"0F",x"49",x"83",
x"CD",x"A4",x"09",x"CD",x"47",x"15",x"C1",x"E1",x"CD",x"A4",x"09",x"EB",x"CD",x"B4",
x"09",x"CD",x"41",x"15",x"C3",x"A0",x"08",x"CD",x"55",x"09",x"FC",x"E2",x"13",x"FC",
x"82",x"09",x"3A",x"24",x"41",x"FE",x"81",x"38",x"0C",x"01",x"00",x"81",x"51",x"59",
x"CD",x"A2",x"08",x"21",x"10",x"07",x"E5",x"21",x"E3",x"15",x"CD",x"9A",x"14",x"21",
x"8B",x"15",x"C9",x"09",x"4A",x"D7",x"3B",x"78",x"02",x"6E",x"84",x"7B",x"FE",x"C1",
x"2F",x"7C",x"74",x"31",x"9A",x"7D",x"84",x"3D",x"5A",x"7D",x"C8",x"7F",x"91",x"7E",
x"E4",x"BB",x"4C",x"7E",x"6C",x"AA",x"AA",x"7F",x"00",x"00",x"00",x"81",x"8A",x"09",
x"37",x"0B",x"77",x"09",x"D4",x"27",x"EF",x"2A",x"F5",x"27",x"E7",x"13",x"C9",x"14",
x"09",x"08",x"39",x"14",x"41",x"15",x"47",x"15",x"A8",x"15",x"BD",x"15",x"AA",x"2C",
x"52",x"41",x"58",x"41",x"5E",x"41",x"61",x"41",x"64",x"41",x"67",x"41",x"6A",x"41",
x"6D",x"41",x"70",x"41",x"7F",x"0A",x"B1",x"0A",x"DB",x"0A",x"26",x"0B",x"03",x"2A",
x"36",x"28",x"C5",x"2A",x"0F",x"2A",x"1F",x"2A",x"61",x"2A",x"91",x"2A",x"9A",x"2A",
x"C5",x"4E",x"44",x"C6",x"4F",x"52",x"D2",x"45",x"53",x"45",x"54",x"D3",x"45",x"54",
x"C3",x"4C",x"53",x"C3",x"4D",x"44",x"D2",x"41",x"4E",x"44",x"4F",x"4D",x"CE",x"45",
x"58",x"54",x"C4",x"41",x"54",x"41",x"C9",x"4E",x"50",x"55",x"54",x"C4",x"49",x"4D",
x"D2",x"45",x"41",x"44",x"CC",x"45",x"54",x"C7",x"4F",x"54",x"4F",x"D2",x"55",x"4E",
x"C9",x"46",x"D2",x"45",x"53",x"54",x"4F",x"52",x"45",x"C7",x"4F",x"53",x"55",x"42",
x"D2",x"45",x"54",x"55",x"52",x"4E",x"D2",x"45",x"4D",x"D3",x"54",x"4F",x"50",x"C5",
x"4C",x"53",x"45",x"D4",x"52",x"4F",x"4E",x"D4",x"52",x"4F",x"46",x"46",x"C4",x"45",
x"46",x"53",x"54",x"52",x"C4",x"45",x"46",x"49",x"4E",x"54",x"C4",x"45",x"46",x"53",
x"4E",x"47",x"C4",x"45",x"46",x"44",x"42",x"4C",x"CC",x"49",x"4E",x"45",x"C5",x"44",
x"49",x"54",x"C5",x"52",x"52",x"4F",x"52",x"D2",x"45",x"53",x"55",x"4D",x"45",x"CF",
x"55",x"54",x"CF",x"4E",x"CF",x"50",x"45",x"4E",x"C6",x"49",x"45",x"4C",x"44",x"C7",
x"45",x"54",x"D0",x"55",x"54",x"C3",x"4C",x"4F",x"53",x"45",x"CC",x"4F",x"41",x"44",
x"CD",x"45",x"52",x"47",x"45",x"CE",x"41",x"4D",x"45",x"CB",x"49",x"4C",x"4C",x"CC",
x"53",x"45",x"54",x"D2",x"53",x"45",x"54",x"D3",x"41",x"56",x"45",x"D3",x"59",x"53",
x"54",x"45",x"4D",x"CC",x"50",x"52",x"49",x"4E",x"54",x"C4",x"45",x"46",x"D0",x"4F",
x"4B",x"45",x"D0",x"52",x"49",x"4E",x"54",x"C3",x"4F",x"4E",x"54",x"CC",x"49",x"53",
x"54",x"CC",x"4C",x"49",x"53",x"54",x"C4",x"45",x"4C",x"45",x"54",x"45",x"C1",x"55",
x"54",x"4F",x"C3",x"4C",x"45",x"41",x"52",x"C3",x"4C",x"4F",x"41",x"44",x"C3",x"53",
x"41",x"56",x"45",x"CE",x"45",x"57",x"D4",x"41",x"42",x"28",x"D4",x"4F",x"C6",x"4E",
x"D5",x"53",x"49",x"4E",x"47",x"D6",x"41",x"52",x"50",x"54",x"52",x"D5",x"53",x"52",
x"C5",x"52",x"4C",x"C5",x"52",x"52",x"D3",x"54",x"52",x"49",x"4E",x"47",x"24",x"C9",
x"4E",x"53",x"54",x"52",x"D0",x"4F",x"49",x"4E",x"54",x"D4",x"49",x"4D",x"45",x"24",
x"CD",x"45",x"4D",x"C9",x"4E",x"4B",x"45",x"59",x"24",x"D4",x"48",x"45",x"4E",x"CE",
x"4F",x"54",x"D3",x"54",x"45",x"50",x"AB",x"AD",x"AA",x"AF",x"DB",x"C1",x"4E",x"44",
x"CF",x"52",x"BE",x"BD",x"BC",x"D3",x"47",x"4E",x"C9",x"4E",x"54",x"C1",x"42",x"53",
x"C6",x"52",x"45",x"C9",x"4E",x"50",x"D0",x"4F",x"53",x"D3",x"51",x"52",x"D2",x"4E",
x"44",x"CC",x"4F",x"47",x"C5",x"58",x"50",x"C3",x"4F",x"53",x"D3",x"49",x"4E",x"D4",
x"41",x"4E",x"C1",x"54",x"4E",x"D0",x"45",x"45",x"4B",x"C3",x"56",x"49",x"C3",x"56",
x"53",x"C3",x"56",x"44",x"C5",x"4F",x"46",x"CC",x"4F",x"43",x"CC",x"4F",x"46",x"CD",
x"4B",x"49",x"24",x"CD",x"4B",x"53",x"24",x"CD",x"4B",x"44",x"24",x"C3",x"49",x"4E",
x"54",x"C3",x"53",x"4E",x"47",x"C3",x"44",x"42",x"4C",x"C6",x"49",x"58",x"CC",x"45",
x"4E",x"D3",x"54",x"52",x"24",x"D6",x"41",x"4C",x"C1",x"53",x"43",x"C3",x"48",x"52",
x"24",x"CC",x"45",x"46",x"54",x"24",x"D2",x"49",x"47",x"48",x"54",x"24",x"CD",x"49",
x"44",x"24",x"A7",x"80",x"AE",x"1D",x"A1",x"1C",x"38",x"01",x"35",x"01",x"C9",x"01",
x"73",x"41",x"D3",x"01",x"B6",x"22",x"05",x"1F",x"9A",x"21",x"08",x"26",x"EF",x"21",
x"21",x"1F",x"C2",x"1E",x"A3",x"1E",x"39",x"20",x"91",x"1D",x"B1",x"1E",x"DE",x"1E",
x"07",x"1F",x"A9",x"1D",x"07",x"1F",x"F7",x"1D",x"F8",x"1D",x"00",x"1E",x"03",x"1E",
x"06",x"1E",x"09",x"1E",x"A3",x"41",x"60",x"2E",x"F4",x"1F",x"AF",x"1F",x"FB",x"2A",
x"6C",x"1F",x"79",x"41",x"7C",x"41",x"7F",x"41",x"82",x"41",x"85",x"41",x"88",x"41",
x"8B",x"41",x"8E",x"41",x"91",x"41",x"97",x"41",x"9A",x"41",x"A0",x"41",x"B2",x"02",
x"67",x"20",x"5B",x"41",x"B1",x"2C",x"6F",x"20",x"E4",x"1D",x"2E",x"2B",x"29",x"2B",
x"C6",x"2B",x"08",x"20",x"7A",x"1E",x"1F",x"2C",x"F5",x"2B",x"49",x"1B",x"79",x"79",
x"7C",x"7C",x"7F",x"50",x"46",x"DB",x"0A",x"00",x"00",x"7F",x"0A",x"F4",x"0A",x"B1",
x"0A",x"77",x"0C",x"70",x"0C",x"A1",x"0D",x"E5",x"0D",x"78",x"0A",x"16",x"07",x"13",
x"07",x"47",x"08",x"A2",x"08",x"0C",x"0A",x"D2",x"0B",x"C7",x"0B",x"F2",x"0B",x"90",
x"24",x"39",x"0A",x"4E",x"46",x"53",x"4E",x"52",x"47",x"4F",x"44",x"46",x"43",x"4F",
x"56",x"4F",x"4D",x"55",x"4C",x"42",x"53",x"44",x"44",x"2F",x"30",x"49",x"44",x"54",
x"4D",x"4F",x"53",x"4C",x"53",x"53",x"54",x"43",x"4E",x"4E",x"52",x"52",x"57",x"55",
x"45",x"4D",x"4F",x"46",x"44",x"53",x"4E",x"D6",x"00",x"6F",x"7C",x"DE",x"00",x"67",
x"78",x"DE",x"00",x"47",x"3E",x"00",x"C9",x"4A",x"1E",x"40",x"E6",x"4D",x"DB",x"00",
x"C9",x"D3",x"00",x"C9",x"00",x"00",x"00",x"00",x"40",x"30",x"00",x"4C",x"43",x"FE",
x"FF",x"E9",x"42",x"20",x"45",x"72",x"72",x"6F",x"72",x"00",x"20",x"69",x"6E",x"20",
x"00",x"52",x"45",x"41",x"44",x"59",x"0D",x"00",x"42",x"72",x"65",x"61",x"6B",x"00",
x"21",x"04",x"00",x"39",x"7E",x"23",x"FE",x"81",x"C0",x"4E",x"23",x"46",x"23",x"E5",
x"69",x"60",x"7A",x"B3",x"EB",x"28",x"02",x"EB",x"DF",x"01",x"0E",x"00",x"E1",x"C8",
x"09",x"18",x"E5",x"CD",x"6C",x"19",x"C5",x"E3",x"C1",x"DF",x"7E",x"02",x"C8",x"0B",
x"2B",x"18",x"F8",x"E5",x"2A",x"FD",x"40",x"06",x"00",x"09",x"09",x"3E",x"E5",x"3E",
x"C6",x"95",x"6F",x"3E",x"FF",x"9C",x"38",x"04",x"67",x"39",x"E1",x"D8",x"1E",x"0C",
x"18",x"24",x"2A",x"A2",x"40",x"7C",x"A5",x"3C",x"28",x"08",x"3A",x"F2",x"40",x"B7",
x"1E",x"22",x"20",x"14",x"C3",x"C1",x"1D",x"2A",x"DA",x"40",x"22",x"A2",x"40",x"1E",
x"02",x"01",x"1E",x"14",x"01",x"1E",x"00",x"01",x"1E",x"24",x"2A",x"A2",x"40",x"22",
x"EA",x"40",x"22",x"EC",x"40",x"01",x"B4",x"19",x"2A",x"E8",x"40",x"C3",x"9A",x"1B",
x"C1",x"7B",x"4B",x"32",x"9A",x"40",x"2A",x"E6",x"40",x"22",x"EE",x"40",x"EB",x"2A",
x"EA",x"40",x"7C",x"A5",x"3C",x"28",x"07",x"22",x"F5",x"40",x"EB",x"22",x"F7",x"40",
x"2A",x"F0",x"40",x"7C",x"B5",x"EB",x"21",x"F2",x"40",x"28",x"08",x"A6",x"20",x"05",
x"35",x"EB",x"C3",x"36",x"1D",x"AF",x"77",x"59",x"CD",x"F9",x"20",x"21",x"C9",x"18",
x"CD",x"A6",x"41",x"57",x"3E",x"3F",x"CD",x"2A",x"03",x"19",x"7E",x"CD",x"2A",x"03",
x"D7",x"CD",x"2A",x"03",x"21",x"1D",x"19",x"E5",x"2A",x"EA",x"40",x"E3",x"CD",x"A7",
x"28",x"E1",x"11",x"FE",x"FF",x"DF",x"CA",x"74",x"06",x"7C",x"A5",x"3C",x"C4",x"A7",
x"0F",x"3E",x"C1",x"CD",x"8B",x"03",x"CD",x"AC",x"41",x"CD",x"F8",x"01",x"CD",x"F9",
x"20",x"21",x"29",x"19",x"CD",x"A7",x"28",x"3A",x"9A",x"40",x"D6",x"02",x"CC",x"53",
x"2E",x"21",x"FF",x"FF",x"22",x"A2",x"40",x"3A",x"E1",x"40",x"B7",x"28",x"37",x"2A",
x"E2",x"40",x"E5",x"CD",x"AF",x"0F",x"D1",x"D5",x"CD",x"2C",x"1B",x"3E",x"2A",x"38",
x"02",x"3E",x"20",x"CD",x"2A",x"03",x"CD",x"61",x"03",x"D1",x"30",x"06",x"AF",x"32",
x"E1",x"40",x"18",x"B9",x"2A",x"E4",x"40",x"19",x"38",x"F4",x"D5",x"11",x"F9",x"FF",
x"DF",x"D1",x"30",x"EC",x"22",x"E2",x"40",x"F6",x"FF",x"C3",x"EB",x"2F",x"3E",x"3E",
x"CD",x"2A",x"03",x"CD",x"61",x"03",x"DA",x"33",x"1A",x"D7",x"3C",x"3D",x"CA",x"33",
x"1A",x"F5",x"CD",x"5A",x"1E",x"2B",x"7E",x"FE",x"20",x"28",x"FA",x"23",x"7E",x"FE",
x"20",x"CC",x"C9",x"09",x"D5",x"CD",x"C0",x"1B",x"D1",x"F1",x"22",x"E6",x"40",x"CD",
x"B2",x"41",x"D2",x"5A",x"1D",x"D5",x"C5",x"AF",x"32",x"DD",x"40",x"D7",x"B7",x"F5",
x"EB",x"22",x"EC",x"40",x"EB",x"CD",x"2C",x"1B",x"C5",x"DC",x"E4",x"2B",x"D1",x"F1",
x"D5",x"28",x"27",x"D1",x"2A",x"F9",x"40",x"E3",x"C1",x"09",x"E5",x"CD",x"55",x"19",
x"E1",x"22",x"F9",x"40",x"EB",x"74",x"D1",x"E5",x"23",x"23",x"73",x"23",x"72",x"23",
x"EB",x"2A",x"A7",x"40",x"EB",x"1B",x"1B",x"1A",x"77",x"23",x"13",x"B7",x"20",x"F9",
x"D1",x"CD",x"FC",x"1A",x"CD",x"B5",x"41",x"CD",x"5D",x"1B",x"CD",x"B8",x"41",x"C3",
x"33",x"1A",x"2A",x"A4",x"40",x"EB",x"62",x"6B",x"7E",x"23",x"B6",x"C8",x"23",x"23",
x"23",x"AF",x"BE",x"23",x"20",x"FC",x"EB",x"73",x"23",x"72",x"18",x"EC",x"11",x"00",
x"00",x"D5",x"28",x"09",x"D1",x"CD",x"4F",x"1E",x"D5",x"28",x"0B",x"CF",x"CE",x"11",
x"FA",x"FF",x"C4",x"4F",x"1E",x"C2",x"97",x"19",x"EB",x"D1",x"E3",x"E5",x"2A",x"A4",
x"40",x"44",x"4D",x"7E",x"23",x"B6",x"2B",x"C8",x"23",x"23",x"7E",x"23",x"66",x"6F",
x"DF",x"60",x"69",x"7E",x"23",x"66",x"6F",x"3F",x"C8",x"3F",x"D0",x"18",x"E6",x"C0",
x"CD",x"C9",x"01",x"2A",x"A4",x"40",x"CD",x"F8",x"1D",x"32",x"E1",x"40",x"77",x"23",
x"77",x"23",x"22",x"F9",x"40",x"2A",x"A4",x"40",x"2B",x"22",x"DF",x"40",x"06",x"1A",
x"21",x"01",x"41",x"36",x"04",x"23",x"10",x"FB",x"AF",x"32",x"F2",x"40",x"6F",x"67",
x"22",x"F0",x"40",x"22",x"F7",x"40",x"2A",x"B1",x"40",x"22",x"D6",x"40",x"CD",x"91",
x"1D",x"2A",x"F9",x"40",x"22",x"FB",x"40",x"22",x"FD",x"40",x"CD",x"BB",x"41",x"C1",
x"2A",x"A0",x"40",x"2B",x"2B",x"22",x"E8",x"40",x"23",x"23",x"F9",x"21",x"B5",x"40",
x"22",x"B3",x"40",x"CD",x"8B",x"03",x"CD",x"69",x"21",x"AF",x"67",x"6F",x"32",x"DC",
x"40",x"E5",x"C5",x"2A",x"DF",x"40",x"C9",x"3E",x"3F",x"CD",x"2A",x"03",x"3E",x"20",
x"CD",x"2A",x"03",x"C3",x"61",x"03",x"AF",x"32",x"B0",x"40",x"4F",x"EB",x"2A",x"A7",
x"40",x"2B",x"2B",x"EB",x"7E",x"FE",x"20",x"CA",x"5B",x"1C",x"47",x"FE",x"22",x"CA",
x"77",x"1C",x"B7",x"CA",x"7D",x"1C",x"3A",x"B0",x"40",x"B7",x"7E",x"C2",x"5B",x"1C",
x"FE",x"3F",x"3E",x"B2",x"CA",x"5B",x"1C",x"7E",x"FE",x"30",x"38",x"05",x"FE",x"3C",
x"DA",x"5B",x"1C",x"D5",x"11",x"4F",x"16",x"C5",x"01",x"3D",x"1C",x"C5",x"06",x"7F",
x"7E",x"FE",x"61",x"38",x"07",x"FE",x"7B",x"30",x"03",x"E6",x"5F",x"77",x"4E",x"EB",
x"23",x"B6",x"F2",x"0E",x"1C",x"04",x"7E",x"E6",x"7F",x"C8",x"B9",x"20",x"F3",x"EB",
x"E5",x"13",x"1A",x"B7",x"FA",x"39",x"1C",x"4F",x"78",x"FE",x"8D",x"20",x"02",x"D7",
x"2B",x"23",x"7E",x"FE",x"61",x"38",x"02",x"E6",x"5F",x"B9",x"28",x"E7",x"E1",x"18",
x"D3",x"48",x"F1",x"EB",x"C9",x"EB",x"79",x"C1",x"D1",x"EB",x"FE",x"95",x"36",x"3A",
x"20",x"02",x"0C",x"23",x"FE",x"FB",x"20",x"0C",x"36",x"3A",x"23",x"06",x"93",x"70",
x"23",x"EB",x"0C",x"0C",x"18",x"1D",x"EB",x"23",x"12",x"13",x"0C",x"D6",x"3A",x"28",
x"04",x"FE",x"4E",x"20",x"03",x"32",x"B0",x"40",x"D6",x"59",x"C2",x"CC",x"1B",x"47",
x"7E",x"B7",x"28",x"09",x"B8",x"28",x"E4",x"23",x"12",x"0C",x"13",x"18",x"F3",x"21",
x"05",x"00",x"44",x"09",x"44",x"4D",x"2A",x"A7",x"40",x"2B",x"2B",x"2B",x"12",x"13",
x"12",x"13",x"12",x"C9",x"7C",x"92",x"C0",x"7D",x"93",x"C9",x"7E",x"E3",x"BE",x"23",
x"E3",x"CA",x"78",x"1D",x"C3",x"97",x"19",x"3E",x"64",x"32",x"DC",x"40",x"CD",x"21",
x"1F",x"E3",x"CD",x"36",x"19",x"D1",x"20",x"05",x"09",x"F9",x"22",x"E8",x"40",x"EB",
x"0E",x"08",x"CD",x"63",x"19",x"E5",x"CD",x"05",x"1F",x"E3",x"E5",x"2A",x"A2",x"40",
x"E3",x"CF",x"BD",x"E7",x"CA",x"F6",x"0A",x"D2",x"F6",x"0A",x"F5",x"CD",x"37",x"23",
x"F1",x"E5",x"F2",x"EC",x"1C",x"CD",x"7F",x"0A",x"E3",x"11",x"01",x"00",x"7E",x"FE",
x"CC",x"CC",x"01",x"2B",x"D5",x"E5",x"EB",x"CD",x"9E",x"09",x"18",x"22",x"CD",x"B1",
x"0A",x"CD",x"BF",x"09",x"E1",x"C5",x"D5",x"01",x"00",x"81",x"51",x"5A",x"7E",x"FE",
x"CC",x"3E",x"01",x"20",x"0E",x"CD",x"38",x"23",x"E5",x"CD",x"B1",x"0A",x"CD",x"BF",
x"09",x"CD",x"55",x"09",x"E1",x"C5",x"D5",x"4F",x"E7",x"47",x"C5",x"E5",x"2A",x"DF",
x"40",x"E3",x"06",x"81",x"C5",x"33",x"CD",x"58",x"03",x"B7",x"C4",x"A0",x"1D",x"22",
x"E6",x"40",x"ED",x"73",x"E8",x"40",x"7E",x"FE",x"3A",x"28",x"29",x"B7",x"C2",x"97",
x"19",x"23",x"7E",x"23",x"B6",x"CA",x"7E",x"19",x"23",x"5E",x"23",x"56",x"EB",x"22",
x"A2",x"40",x"3A",x"1B",x"41",x"B7",x"28",x"0F",x"D5",x"3E",x"3C",x"CD",x"2A",x"03",
x"CD",x"AF",x"0F",x"3E",x"3E",x"CD",x"2A",x"03",x"D1",x"EB",x"D7",x"11",x"1E",x"1D",
x"D5",x"C8",x"D6",x"80",x"DA",x"21",x"1F",x"FE",x"3C",x"D2",x"E7",x"2A",x"07",x"4F",
x"06",x"00",x"EB",x"21",x"22",x"18",x"09",x"4E",x"23",x"46",x"C5",x"EB",x"23",x"7E",
x"FE",x"3A",x"D0",x"FE",x"20",x"CA",x"78",x"1D",x"FE",x"0B",x"30",x"05",x"FE",x"09",
x"D2",x"78",x"1D",x"FE",x"30",x"3F",x"3C",x"3D",x"C9",x"EB",x"2A",x"A4",x"40",x"2B",
x"22",x"FF",x"40",x"EB",x"C9",x"CD",x"58",x"03",x"B7",x"C8",x"FE",x"60",x"CC",x"84",
x"03",x"32",x"99",x"40",x"3D",x"C0",x"3C",x"C3",x"B4",x"1D",x"C0",x"F5",x"CC",x"BB",
x"41",x"F1",x"22",x"E6",x"40",x"21",x"B5",x"40",x"22",x"B3",x"40",x"21",x"F6",x"FF",
x"C1",x"2A",x"A2",x"40",x"E5",x"F5",x"7D",x"A4",x"3C",x"28",x"09",x"22",x"F5",x"40",
x"2A",x"E6",x"40",x"22",x"F7",x"40",x"CD",x"8B",x"03",x"CD",x"F9",x"20",x"F1",x"21",
x"30",x"19",x"C2",x"06",x"1A",x"C3",x"18",x"1A",x"2A",x"F7",x"40",x"7C",x"B5",x"1E",
x"20",x"CA",x"A2",x"19",x"EB",x"2A",x"F5",x"40",x"22",x"A2",x"40",x"EB",x"C9",x"3E",
x"AF",x"32",x"1B",x"41",x"C9",x"F1",x"E1",x"C9",x"1E",x"03",x"01",x"1E",x"02",x"01",
x"1E",x"04",x"01",x"1E",x"08",x"CD",x"3D",x"1E",x"01",x"97",x"19",x"C5",x"D8",x"D6",
x"41",x"4F",x"47",x"D7",x"FE",x"CE",x"20",x"09",x"D7",x"CD",x"3D",x"1E",x"D8",x"D6",
x"41",x"47",x"D7",x"78",x"91",x"D8",x"3C",x"E3",x"21",x"01",x"41",x"06",x"00",x"09",
x"73",x"23",x"3D",x"20",x"FB",x"E1",x"7E",x"FE",x"2C",x"C0",x"D7",x"18",x"CE",x"7E",
x"FE",x"41",x"D8",x"FE",x"5B",x"3F",x"C9",x"D7",x"CD",x"02",x"2B",x"F0",x"1E",x"08",
x"C3",x"A2",x"19",x"7E",x"FE",x"2E",x"EB",x"2A",x"EC",x"40",x"EB",x"CA",x"78",x"1D",
x"2B",x"11",x"00",x"00",x"D7",x"D0",x"E5",x"F5",x"21",x"98",x"19",x"DF",x"DA",x"97",
x"19",x"62",x"6B",x"19",x"29",x"19",x"29",x"F1",x"D6",x"30",x"5F",x"16",x"00",x"19",
x"EB",x"E1",x"18",x"E4",x"CA",x"61",x"1B",x"CD",x"46",x"1E",x"2B",x"D7",x"C0",x"E5",
x"2A",x"B1",x"40",x"7D",x"93",x"5F",x"7C",x"9A",x"57",x"DA",x"7A",x"19",x"2A",x"F9",
x"40",x"01",x"28",x"00",x"09",x"DF",x"D2",x"7A",x"19",x"EB",x"22",x"A0",x"40",x"E1",
x"C3",x"61",x"1B",x"CA",x"5D",x"1B",x"CD",x"C7",x"41",x"CD",x"61",x"1B",x"01",x"1E",
x"1D",x"18",x"10",x"0E",x"03",x"CD",x"63",x"19",x"C1",x"E5",x"E5",x"2A",x"A2",x"40",
x"E3",x"3E",x"91",x"F5",x"33",x"C5",x"CD",x"5A",x"1E",x"CD",x"07",x"1F",x"E5",x"2A",
x"A2",x"40",x"DF",x"E1",x"23",x"DC",x"2F",x"1B",x"D4",x"2C",x"1B",x"60",x"69",x"2B",
x"D8",x"1E",x"0E",x"C3",x"A2",x"19",x"C0",x"16",x"FF",x"CD",x"36",x"19",x"F9",x"22",
x"E8",x"40",x"FE",x"91",x"1E",x"04",x"C2",x"A2",x"19",x"E1",x"22",x"A2",x"40",x"23",
x"7C",x"B5",x"20",x"07",x"3A",x"DD",x"40",x"B7",x"C2",x"18",x"1A",x"21",x"1E",x"1D",
x"E3",x"3E",x"E1",x"01",x"3A",x"0E",x"00",x"06",x"00",x"79",x"48",x"47",x"7E",x"B7",
x"C8",x"B8",x"C8",x"23",x"FE",x"22",x"28",x"F3",x"D6",x"8F",x"20",x"F2",x"B8",x"8A",
x"57",x"18",x"ED",x"CD",x"0D",x"26",x"CF",x"D5",x"EB",x"22",x"DF",x"40",x"EB",x"D5",
x"E7",x"F5",x"CD",x"37",x"23",x"F1",x"E3",x"C6",x"03",x"CD",x"19",x"28",x"CD",x"03",
x"0A",x"E5",x"20",x"28",x"2A",x"21",x"41",x"E5",x"23",x"5E",x"23",x"56",x"2A",x"A4",
x"40",x"DF",x"30",x"0E",x"2A",x"A0",x"40",x"DF",x"D1",x"30",x"0F",x"2A",x"F9",x"40",
x"DF",x"30",x"09",x"3E",x"D1",x"CD",x"F5",x"29",x"EB",x"CD",x"43",x"28",x"CD",x"F5",
x"29",x"E3",x"CD",x"D3",x"09",x"D1",x"E1",x"C9",x"FE",x"9E",x"20",x"25",x"D7",x"CF",
x"8D",x"CD",x"5A",x"1E",x"7A",x"B3",x"28",x"09",x"CD",x"2A",x"1B",x"50",x"59",x"E1",
x"D2",x"D9",x"1E",x"EB",x"22",x"F0",x"40",x"EB",x"D8",x"3A",x"F2",x"40",x"B7",x"C8",
x"3A",x"9A",x"40",x"5F",x"C3",x"AB",x"19",x"CD",x"1C",x"2B",x"7E",x"47",x"FE",x"91",
x"28",x"03",x"CF",x"8D",x"2B",x"4B",x"0D",x"78",x"CA",x"60",x"1D",x"CD",x"5B",x"1E",
x"FE",x"2C",x"C0",x"18",x"F3",x"11",x"F2",x"40",x"1A",x"B7",x"CA",x"A0",x"19",x"3C",
x"32",x"9A",x"40",x"12",x"7E",x"FE",x"87",x"28",x"0C",x"CD",x"5A",x"1E",x"C0",x"7A",
x"B3",x"C2",x"C5",x"1E",x"3C",x"18",x"02",x"D7",x"C0",x"2A",x"EE",x"40",x"EB",x"2A",
x"EA",x"40",x"22",x"A2",x"40",x"EB",x"C0",x"7E",x"B7",x"20",x"04",x"23",x"23",x"23",
x"23",x"23",x"7A",x"A3",x"3C",x"C2",x"05",x"1F",x"3A",x"DD",x"40",x"3D",x"CA",x"BE",
x"1D",x"C3",x"05",x"1F",x"CD",x"1C",x"2B",x"C0",x"B7",x"CA",x"4A",x"1E",x"3D",x"87",
x"5F",x"FE",x"2D",x"38",x"02",x"1E",x"26",x"C3",x"A2",x"19",x"11",x"0A",x"00",x"D5",
x"28",x"17",x"CD",x"4F",x"1E",x"EB",x"E3",x"28",x"11",x"EB",x"CF",x"2C",x"EB",x"2A",
x"E4",x"40",x"EB",x"28",x"06",x"CD",x"5A",x"1E",x"C2",x"97",x"19",x"EB",x"7C",x"B5",
x"CA",x"4A",x"1E",x"22",x"E4",x"40",x"32",x"E1",x"40",x"E1",x"22",x"E2",x"40",x"C1",
x"C3",x"33",x"1A",x"CD",x"37",x"23",x"7E",x"FE",x"2C",x"CC",x"78",x"1D",x"FE",x"CA",
x"CC",x"78",x"1D",x"2B",x"E5",x"CD",x"94",x"09",x"E1",x"28",x"07",x"D7",x"DA",x"C2",
x"1E",x"C3",x"5F",x"1D",x"16",x"01",x"CD",x"05",x"1F",x"B7",x"C8",x"D7",x"FE",x"95",
x"20",x"F6",x"15",x"20",x"F3",x"18",x"E8",x"3E",x"01",x"32",x"9C",x"40",x"C3",x"9B",
x"20",x"CD",x"CA",x"41",x"FE",x"40",x"20",x"19",x"CD",x"01",x"2B",x"FE",x"04",x"D2",
x"4A",x"1E",x"E5",x"21",x"00",x"3C",x"19",x"22",x"20",x"40",x"7B",x"E6",x"3F",x"32",
x"A6",x"40",x"E1",x"CF",x"2C",x"FE",x"23",x"20",x"08",x"CD",x"84",x"02",x"3E",x"80",
x"32",x"9C",x"40",x"2B",x"D7",x"CC",x"FE",x"20",x"CA",x"69",x"21",x"FE",x"BF",x"CA",
x"BD",x"2C",x"FE",x"BC",x"CA",x"37",x"21",x"E5",x"FE",x"2C",x"CA",x"08",x"21",x"FE",
x"3B",x"CA",x"64",x"21",x"C1",x"CD",x"37",x"23",x"E5",x"E7",x"28",x"32",x"CD",x"BD",
x"0F",x"CD",x"65",x"28",x"CD",x"CD",x"41",x"2A",x"21",x"41",x"3A",x"9C",x"40",x"B7",
x"FA",x"E9",x"20",x"28",x"08",x"3A",x"9B",x"40",x"86",x"FE",x"84",x"18",x"09",x"3A",
x"9D",x"40",x"47",x"3A",x"A6",x"40",x"86",x"B8",x"D4",x"FE",x"20",x"CD",x"AA",x"28",
x"3E",x"20",x"CD",x"2A",x"03",x"B7",x"CC",x"AA",x"28",x"E1",x"C3",x"9B",x"20",x"3A",
x"A6",x"40",x"B7",x"C8",x"3E",x"0D",x"CD",x"2A",x"03",x"CD",x"D0",x"41",x"AF",x"C9",
x"CD",x"D3",x"41",x"3A",x"9C",x"40",x"B7",x"F2",x"19",x"21",x"3E",x"2C",x"CD",x"2A",
x"03",x"18",x"4B",x"28",x"08",x"3A",x"9B",x"40",x"FE",x"70",x"C3",x"2B",x"21",x"3A",
x"9E",x"40",x"47",x"3A",x"A6",x"40",x"B8",x"D4",x"FE",x"20",x"30",x"34",x"D6",x"10",
x"30",x"FC",x"2F",x"18",x"23",x"CD",x"1B",x"2B",x"E6",x"3F",x"5F",x"CF",x"29",x"2B",
x"E5",x"CD",x"D3",x"41",x"3A",x"9C",x"40",x"B7",x"FA",x"4A",x"1E",x"CA",x"53",x"21",
x"3A",x"9B",x"40",x"18",x"03",x"3A",x"A6",x"40",x"2F",x"83",x"30",x"0A",x"3C",x"47",
x"3E",x"20",x"CD",x"2A",x"03",x"05",x"20",x"FA",x"E1",x"D7",x"C3",x"A0",x"20",x"3A",
x"9C",x"40",x"B7",x"FC",x"F8",x"01",x"AF",x"32",x"9C",x"40",x"CD",x"BE",x"41",x"C9",
x"3F",x"52",x"45",x"44",x"4F",x"0D",x"00",x"3A",x"DE",x"40",x"B7",x"C2",x"91",x"19",
x"3A",x"A9",x"40",x"B7",x"1E",x"2A",x"CA",x"A2",x"19",x"C1",x"21",x"78",x"21",x"CD",
x"A7",x"28",x"2A",x"E6",x"40",x"C9",x"CD",x"28",x"28",x"7E",x"CD",x"D6",x"41",x"D6",
x"23",x"32",x"A9",x"40",x"7E",x"20",x"20",x"CD",x"93",x"02",x"E5",x"06",x"FA",x"2A",
x"A7",x"40",x"CD",x"35",x"02",x"77",x"23",x"FE",x"0D",x"28",x"02",x"10",x"F5",x"2B",
x"36",x"00",x"CD",x"F8",x"01",x"2A",x"A7",x"40",x"2B",x"18",x"22",x"01",x"DB",x"21",
x"C5",x"FE",x"22",x"C0",x"CD",x"66",x"28",x"CF",x"3B",x"E5",x"CD",x"AA",x"28",x"E1",
x"C9",x"E5",x"CD",x"B3",x"1B",x"C1",x"DA",x"BE",x"1D",x"23",x"7E",x"B7",x"2B",x"C5",
x"CA",x"04",x"1F",x"36",x"2C",x"18",x"05",x"E5",x"2A",x"FF",x"40",x"F6",x"AF",x"32",
x"DE",x"40",x"E3",x"18",x"02",x"CF",x"2C",x"CD",x"0D",x"26",x"E3",x"D5",x"7E",x"FE",
x"2C",x"28",x"26",x"3A",x"DE",x"40",x"B7",x"C2",x"96",x"22",x"3A",x"A9",x"40",x"B7",
x"1E",x"06",x"CA",x"A2",x"19",x"3E",x"3F",x"CD",x"2A",x"03",x"CD",x"B3",x"1B",x"D1",
x"C1",x"DA",x"BE",x"1D",x"23",x"7E",x"B7",x"2B",x"C5",x"CA",x"04",x"1F",x"D5",x"CD",
x"DC",x"41",x"E7",x"F5",x"20",x"19",x"D7",x"57",x"47",x"FE",x"22",x"28",x"05",x"16",
x"3A",x"06",x"2C",x"2B",x"CD",x"69",x"28",x"F1",x"EB",x"21",x"5A",x"22",x"E3",x"D5",
x"C3",x"33",x"1F",x"D7",x"F1",x"F5",x"01",x"43",x"22",x"C5",x"DA",x"6C",x"0E",x"D2",
x"65",x"0E",x"2B",x"D7",x"28",x"05",x"FE",x"2C",x"C2",x"7F",x"21",x"E3",x"2B",x"D7",
x"C2",x"FB",x"21",x"D1",x"00",x"00",x"00",x"00",x"00",x"3A",x"DE",x"40",x"B7",x"EB",
x"C2",x"96",x"1D",x"D5",x"CD",x"DF",x"41",x"B6",x"21",x"86",x"22",x"C4",x"A7",x"28",
x"E1",x"C3",x"69",x"21",x"3F",x"45",x"78",x"74",x"72",x"61",x"20",x"69",x"67",x"6E",
x"6F",x"72",x"65",x"64",x"0D",x"00",x"CD",x"05",x"1F",x"B7",x"20",x"12",x"23",x"7E",
x"23",x"B6",x"1E",x"06",x"CA",x"A2",x"19",x"23",x"5E",x"23",x"56",x"EB",x"22",x"DA",
x"40",x"EB",x"D7",x"FE",x"88",x"20",x"E3",x"C3",x"2D",x"22",x"11",x"00",x"00",x"C4",
x"0D",x"26",x"22",x"DF",x"40",x"CD",x"36",x"19",x"C2",x"9D",x"19",x"F9",x"22",x"E8",
x"40",x"D5",x"7E",x"23",x"F5",x"D5",x"7E",x"23",x"B7",x"FA",x"EA",x"22",x"CD",x"B1",
x"09",x"E3",x"E5",x"CD",x"0B",x"07",x"E1",x"CD",x"CB",x"09",x"E1",x"CD",x"C2",x"09",
x"E5",x"CD",x"0C",x"0A",x"18",x"29",x"23",x"23",x"23",x"23",x"4E",x"23",x"46",x"23",
x"E3",x"5E",x"23",x"56",x"E5",x"69",x"60",x"CD",x"D2",x"0B",x"3A",x"AF",x"40",x"FE",
x"04",x"CA",x"B2",x"07",x"EB",x"E1",x"72",x"2B",x"73",x"E1",x"D5",x"5E",x"23",x"56",
x"23",x"E3",x"CD",x"39",x"0A",x"E1",x"C1",x"90",x"CD",x"C2",x"09",x"28",x"09",x"EB",
x"22",x"A2",x"40",x"69",x"60",x"C3",x"1A",x"1D",x"F9",x"22",x"E8",x"40",x"2A",x"DF",
x"40",x"7E",x"FE",x"2C",x"C2",x"1E",x"1D",x"D7",x"CD",x"B9",x"22",x"CF",x"28",x"2B",
x"16",x"00",x"D5",x"0E",x"01",x"CD",x"63",x"19",x"CD",x"9F",x"24",x"22",x"F3",x"40",
x"2A",x"F3",x"40",x"C1",x"7E",x"16",x"00",x"D6",x"D4",x"38",x"13",x"FE",x"03",x"30",
x"0F",x"FE",x"01",x"17",x"AA",x"BA",x"57",x"DA",x"97",x"19",x"22",x"D8",x"40",x"D7",
x"18",x"E9",x"7A",x"B7",x"C2",x"EC",x"23",x"7E",x"22",x"D8",x"40",x"D6",x"CD",x"D8",
x"FE",x"07",x"D0",x"5F",x"3A",x"AF",x"40",x"D6",x"03",x"B3",x"CA",x"8F",x"29",x"21",
x"9A",x"18",x"19",x"78",x"56",x"BA",x"D0",x"C5",x"01",x"46",x"23",x"C5",x"7A",x"FE",
x"7F",x"CA",x"D4",x"23",x"FE",x"51",x"DA",x"E1",x"23",x"21",x"21",x"41",x"B7",x"3A",
x"AF",x"40",x"3D",x"3D",x"3D",x"CA",x"F6",x"0A",x"4E",x"23",x"46",x"C5",x"FA",x"C5",
x"23",x"23",x"4E",x"23",x"46",x"C5",x"F5",x"B7",x"E2",x"C4",x"23",x"F1",x"23",x"38",
x"03",x"21",x"1D",x"41",x"4E",x"23",x"46",x"23",x"C5",x"4E",x"23",x"46",x"C5",x"06",
x"F1",x"C6",x"03",x"4B",x"47",x"C5",x"01",x"06",x"24",x"C5",x"2A",x"D8",x"40",x"C3",
x"3A",x"23",x"CD",x"B1",x"0A",x"CD",x"A4",x"09",x"01",x"F2",x"13",x"16",x"7F",x"18",
x"EC",x"D5",x"CD",x"7F",x"0A",x"D1",x"E5",x"01",x"E9",x"25",x"18",x"E1",x"78",x"FE",
x"64",x"D0",x"C5",x"D5",x"11",x"04",x"64",x"21",x"B8",x"25",x"E5",x"E7",x"C2",x"95",
x"23",x"2A",x"21",x"41",x"E5",x"01",x"8C",x"25",x"18",x"C7",x"C1",x"79",x"32",x"B0",
x"40",x"78",x"FE",x"08",x"28",x"28",x"3A",x"AF",x"40",x"FE",x"08",x"CA",x"60",x"24",
x"57",x"78",x"FE",x"04",x"CA",x"72",x"24",x"7A",x"FE",x"03",x"CA",x"F6",x"0A",x"D2",
x"7C",x"24",x"21",x"BF",x"18",x"06",x"00",x"09",x"09",x"4E",x"23",x"46",x"D1",x"2A",
x"21",x"41",x"C5",x"C9",x"CD",x"DB",x"0A",x"CD",x"FC",x"09",x"E1",x"22",x"1F",x"41",
x"E1",x"22",x"1D",x"41",x"C1",x"D1",x"CD",x"B4",x"09",x"CD",x"DB",x"0A",x"21",x"AB",
x"18",x"3A",x"B0",x"40",x"07",x"C5",x"4F",x"06",x"00",x"09",x"C1",x"7E",x"23",x"66",
x"6F",x"E9",x"C5",x"CD",x"FC",x"09",x"F1",x"32",x"AF",x"40",x"FE",x"04",x"28",x"DA",
x"E1",x"22",x"21",x"41",x"18",x"D9",x"CD",x"B1",x"0A",x"C1",x"D1",x"21",x"B5",x"18",
x"18",x"D5",x"E1",x"CD",x"A4",x"09",x"CD",x"CF",x"0A",x"CD",x"BF",x"09",x"E1",x"22",
x"23",x"41",x"E1",x"22",x"21",x"41",x"18",x"E7",x"E5",x"EB",x"CD",x"CF",x"0A",x"E1",
x"CD",x"A4",x"09",x"CD",x"CF",x"0A",x"C3",x"A0",x"08",x"D7",x"1E",x"28",x"CA",x"A2",
x"19",x"DA",x"6C",x"0E",x"CD",x"3D",x"1E",x"D2",x"40",x"25",x"FE",x"CD",x"28",x"ED",
x"FE",x"2E",x"CA",x"6C",x"0E",x"FE",x"CE",x"CA",x"32",x"25",x"FE",x"22",x"CA",x"66",
x"28",x"FE",x"CB",x"CA",x"C4",x"25",x"FE",x"26",x"CA",x"94",x"41",x"FE",x"C3",x"20",
x"0A",x"D7",x"3A",x"9A",x"40",x"E5",x"CD",x"F8",x"27",x"E1",x"C9",x"FE",x"C2",x"20",
x"0A",x"D7",x"E5",x"2A",x"EA",x"40",x"CD",x"66",x"0C",x"E1",x"C9",x"FE",x"C0",x"20",
x"14",x"D7",x"CF",x"28",x"CD",x"0D",x"26",x"CF",x"29",x"E5",x"EB",x"7C",x"B5",x"CA",
x"4A",x"1E",x"CD",x"9A",x"0A",x"E1",x"C9",x"FE",x"C1",x"CA",x"FE",x"27",x"FE",x"C5",
x"CA",x"9D",x"41",x"FE",x"C8",x"CA",x"C9",x"27",x"FE",x"C7",x"CA",x"76",x"41",x"FE",
x"C6",x"CA",x"32",x"01",x"FE",x"C9",x"CA",x"9D",x"01",x"FE",x"C4",x"CA",x"2F",x"2A",
x"FE",x"BE",x"CA",x"55",x"41",x"D6",x"D7",x"D2",x"4E",x"25",x"CD",x"35",x"23",x"CF",
x"29",x"C9",x"16",x"7D",x"CD",x"3A",x"23",x"2A",x"F3",x"40",x"E5",x"CD",x"7B",x"09",
x"E1",x"C9",x"CD",x"0D",x"26",x"E5",x"EB",x"22",x"21",x"41",x"E7",x"C4",x"F7",x"09",
x"E1",x"C9",x"06",x"00",x"07",x"4F",x"C5",x"D7",x"79",x"FE",x"41",x"38",x"16",x"CD",
x"35",x"23",x"CF",x"2C",x"CD",x"F4",x"0A",x"EB",x"2A",x"21",x"41",x"E3",x"E5",x"EB",
x"CD",x"1C",x"2B",x"EB",x"E3",x"18",x"14",x"CD",x"2C",x"25",x"E3",x"7D",x"FE",x"0C",
x"38",x"07",x"FE",x"1B",x"E5",x"DC",x"B1",x"0A",x"E1",x"11",x"3E",x"25",x"D5",x"01",
x"08",x"16",x"09",x"4E",x"23",x"66",x"69",x"E9",x"CD",x"D7",x"29",x"7E",x"23",x"4E",
x"23",x"46",x"D1",x"C5",x"F5",x"CD",x"DE",x"29",x"D1",x"5E",x"23",x"4E",x"23",x"46",
x"E1",x"7B",x"B2",x"C8",x"7A",x"D6",x"01",x"D8",x"AF",x"BB",x"3C",x"D0",x"15",x"1D",
x"0A",x"BE",x"23",x"03",x"28",x"ED",x"3F",x"C3",x"60",x"09",x"3C",x"8F",x"C1",x"A0",
x"C6",x"FF",x"9F",x"CD",x"8D",x"09",x"18",x"12",x"16",x"5A",x"CD",x"3A",x"23",x"CD",
x"7F",x"0A",x"7D",x"2F",x"6F",x"7C",x"2F",x"67",x"22",x"21",x"41",x"C1",x"C3",x"46",
x"23",x"3A",x"AF",x"40",x"FE",x"08",x"30",x"05",x"D6",x"03",x"B7",x"37",x"C9",x"D6",
x"03",x"B7",x"C9",x"C5",x"CD",x"7F",x"0A",x"F1",x"D1",x"01",x"FA",x"27",x"C5",x"FE",
x"46",x"20",x"06",x"7B",x"B5",x"6F",x"7C",x"B2",x"C9",x"7B",x"A5",x"6F",x"7C",x"A2",
x"C9",x"2B",x"D7",x"C8",x"CF",x"2C",x"01",x"03",x"26",x"C5",x"F6",x"AF",x"32",x"AE",
x"40",x"46",x"CD",x"3D",x"1E",x"DA",x"97",x"19",x"AF",x"4F",x"D7",x"38",x"05",x"CD",
x"3D",x"1E",x"38",x"09",x"4F",x"D7",x"38",x"FD",x"CD",x"3D",x"1E",x"30",x"F8",x"11",
x"52",x"26",x"D5",x"16",x"02",x"FE",x"25",x"C8",x"14",x"FE",x"24",x"C8",x"14",x"FE",
x"21",x"C8",x"16",x"08",x"FE",x"23",x"C8",x"78",x"D6",x"41",x"E6",x"7F",x"5F",x"16",
x"00",x"E5",x"21",x"01",x"41",x"19",x"56",x"E1",x"2B",x"C9",x"7A",x"32",x"AF",x"40",
x"D7",x"3A",x"DC",x"40",x"B7",x"C2",x"64",x"26",x"7E",x"D6",x"28",x"CA",x"E9",x"26",
x"AF",x"32",x"DC",x"40",x"E5",x"D5",x"2A",x"F9",x"40",x"EB",x"2A",x"FB",x"40",x"DF",
x"E1",x"28",x"19",x"1A",x"6F",x"BC",x"13",x"20",x"0B",x"1A",x"B9",x"20",x"07",x"13",
x"1A",x"B8",x"CA",x"CC",x"26",x"3E",x"13",x"13",x"E5",x"26",x"00",x"19",x"18",x"DF",
x"7C",x"E1",x"E3",x"F5",x"D5",x"11",x"F1",x"24",x"DF",x"28",x"36",x"11",x"43",x"25",
x"DF",x"D1",x"28",x"35",x"F1",x"E3",x"E5",x"C5",x"4F",x"06",x"00",x"C5",x"03",x"03",
x"03",x"2A",x"FD",x"40",x"E5",x"09",x"C1",x"E5",x"CD",x"55",x"19",x"E1",x"22",x"FD",
x"40",x"60",x"69",x"22",x"FB",x"40",x"2B",x"36",x"00",x"DF",x"20",x"FA",x"D1",x"73",
x"23",x"D1",x"73",x"23",x"72",x"EB",x"13",x"E1",x"C9",x"57",x"5F",x"F1",x"F1",x"E3",
x"C9",x"32",x"24",x"41",x"C1",x"67",x"6F",x"22",x"21",x"41",x"E7",x"20",x"06",x"21",
x"28",x"19",x"22",x"21",x"41",x"E1",x"C9",x"E5",x"2A",x"AE",x"40",x"E3",x"57",x"D5",
x"C5",x"CD",x"45",x"1E",x"C1",x"F1",x"EB",x"E3",x"E5",x"EB",x"3C",x"57",x"7E",x"FE",
x"2C",x"28",x"EE",x"CF",x"29",x"22",x"F3",x"40",x"E1",x"22",x"AE",x"40",x"D5",x"2A",
x"FB",x"40",x"3E",x"19",x"EB",x"2A",x"FD",x"40",x"EB",x"DF",x"3A",x"AF",x"40",x"28",
x"27",x"BE",x"23",x"20",x"08",x"7E",x"B9",x"23",x"20",x"04",x"7E",x"B8",x"3E",x"23",
x"23",x"5E",x"23",x"56",x"23",x"20",x"E0",x"3A",x"AE",x"40",x"B7",x"1E",x"12",x"C2",
x"A2",x"19",x"F1",x"96",x"CA",x"95",x"27",x"1E",x"10",x"C3",x"A2",x"19",x"77",x"23",
x"5F",x"16",x"00",x"F1",x"71",x"23",x"70",x"23",x"4F",x"CD",x"63",x"19",x"23",x"23",
x"22",x"D8",x"40",x"71",x"23",x"3A",x"AE",x"40",x"17",x"79",x"01",x"0B",x"00",x"30",
x"02",x"C1",x"03",x"71",x"23",x"70",x"23",x"F5",x"CD",x"AA",x"0B",x"F1",x"3D",x"20",
x"ED",x"F5",x"42",x"4B",x"EB",x"19",x"38",x"C7",x"CD",x"6C",x"19",x"22",x"FD",x"40",
x"2B",x"36",x"00",x"DF",x"20",x"FA",x"03",x"57",x"2A",x"D8",x"40",x"5E",x"EB",x"29",
x"09",x"EB",x"2B",x"2B",x"73",x"23",x"72",x"23",x"F1",x"38",x"30",x"47",x"4F",x"7E",
x"23",x"16",x"E1",x"5E",x"23",x"56",x"23",x"E3",x"F5",x"DF",x"D2",x"3D",x"27",x"CD",
x"AA",x"0B",x"19",x"F1",x"3D",x"44",x"4D",x"20",x"EB",x"3A",x"AF",x"40",x"44",x"4D",
x"29",x"D6",x"04",x"38",x"04",x"29",x"28",x"06",x"29",x"B7",x"E2",x"C2",x"27",x"09",
x"C1",x"09",x"EB",x"2A",x"F3",x"40",x"C9",x"AF",x"E5",x"32",x"AF",x"40",x"CD",x"D4",
x"27",x"E1",x"D7",x"C9",x"2A",x"FD",x"40",x"EB",x"21",x"00",x"00",x"39",x"E7",x"20",
x"0D",x"CD",x"DA",x"29",x"CD",x"E6",x"28",x"2A",x"A0",x"40",x"EB",x"2A",x"D6",x"40",
x"7D",x"93",x"6F",x"7C",x"9A",x"67",x"C3",x"66",x"0C",x"3A",x"A6",x"40",x"6F",x"AF",
x"67",x"C3",x"9A",x"0A",x"CD",x"A9",x"41",x"D7",x"CD",x"2C",x"25",x"E5",x"21",x"90",
x"08",x"E5",x"3A",x"AF",x"40",x"F5",x"FE",x"03",x"CC",x"DA",x"29",x"F1",x"EB",x"2A",
x"8E",x"40",x"E9",x"E5",x"E6",x"07",x"21",x"A1",x"18",x"4F",x"06",x"00",x"09",x"CD",
x"86",x"25",x"E1",x"C9",x"E5",x"2A",x"A2",x"40",x"23",x"7C",x"B5",x"E1",x"C0",x"1E",
x"16",x"C3",x"A2",x"19",x"CD",x"BD",x"0F",x"CD",x"65",x"28",x"CD",x"DA",x"29",x"01",
x"2B",x"2A",x"C5",x"7E",x"23",x"E5",x"CD",x"BF",x"28",x"E1",x"4E",x"23",x"46",x"CD",
x"5A",x"28",x"E5",x"6F",x"CD",x"CE",x"29",x"D1",x"C9",x"CD",x"BF",x"28",x"21",x"D3",
x"40",x"E5",x"77",x"23",x"73",x"23",x"72",x"E1",x"C9",x"2B",x"06",x"22",x"50",x"E5",
x"0E",x"FF",x"23",x"7E",x"0C",x"B7",x"28",x"06",x"BA",x"28",x"03",x"B8",x"20",x"F4",
x"FE",x"22",x"CC",x"78",x"1D",x"E3",x"23",x"EB",x"79",x"CD",x"5A",x"28",x"11",x"D3",
x"40",x"3E",x"D5",x"2A",x"B3",x"40",x"22",x"21",x"41",x"3E",x"03",x"32",x"AF",x"40",
x"CD",x"D3",x"09",x"11",x"D6",x"40",x"DF",x"22",x"B3",x"40",x"E1",x"7E",x"C0",x"1E",
x"1E",x"C3",x"A2",x"19",x"23",x"CD",x"65",x"28",x"CD",x"DA",x"29",x"CD",x"C4",x"09",
x"14",x"15",x"C8",x"0A",x"CD",x"2A",x"03",x"FE",x"0D",x"CC",x"03",x"21",x"03",x"18",
x"F2",x"B7",x"0E",x"F1",x"F5",x"2A",x"A0",x"40",x"EB",x"2A",x"D6",x"40",x"2F",x"4F",
x"06",x"FF",x"09",x"23",x"DF",x"38",x"07",x"22",x"D6",x"40",x"23",x"EB",x"F1",x"C9",
x"F1",x"1E",x"1A",x"CA",x"A2",x"19",x"BF",x"F5",x"01",x"C1",x"28",x"C5",x"2A",x"B1",
x"40",x"22",x"D6",x"40",x"21",x"00",x"00",x"E5",x"2A",x"A0",x"40",x"E5",x"21",x"B5",
x"40",x"EB",x"2A",x"B3",x"40",x"EB",x"DF",x"01",x"F7",x"28",x"C2",x"4A",x"29",x"2A",
x"F9",x"40",x"EB",x"2A",x"FB",x"40",x"EB",x"DF",x"28",x"13",x"7E",x"23",x"23",x"23",
x"FE",x"03",x"20",x"04",x"CD",x"4B",x"29",x"AF",x"5F",x"16",x"00",x"19",x"18",x"E6",
x"C1",x"EB",x"2A",x"FD",x"40",x"EB",x"DF",x"CA",x"6B",x"29",x"7E",x"23",x"CD",x"C2",
x"09",x"E5",x"09",x"FE",x"03",x"20",x"EB",x"22",x"D8",x"40",x"E1",x"4E",x"06",x"00",
x"09",x"09",x"23",x"EB",x"2A",x"D8",x"40",x"EB",x"DF",x"28",x"DA",x"01",x"3F",x"29",
x"C5",x"AF",x"B6",x"23",x"5E",x"23",x"56",x"23",x"C8",x"44",x"4D",x"2A",x"D6",x"40",
x"DF",x"60",x"69",x"D8",x"E1",x"E3",x"DF",x"E3",x"E5",x"60",x"69",x"D0",x"C1",x"F1",
x"F1",x"E5",x"D5",x"C5",x"C9",x"D1",x"E1",x"7D",x"B4",x"C8",x"2B",x"46",x"2B",x"4E",
x"E5",x"2B",x"6E",x"26",x"00",x"09",x"50",x"59",x"2B",x"44",x"4D",x"2A",x"D6",x"40",
x"CD",x"58",x"19",x"E1",x"71",x"23",x"70",x"69",x"60",x"2B",x"C3",x"E9",x"28",x"C5",
x"E5",x"2A",x"21",x"41",x"E3",x"CD",x"9F",x"24",x"E3",x"CD",x"F4",x"0A",x"7E",x"E5",
x"2A",x"21",x"41",x"E5",x"86",x"1E",x"1C",x"DA",x"A2",x"19",x"CD",x"57",x"28",x"D1",
x"CD",x"DE",x"29",x"E3",x"CD",x"DD",x"29",x"E5",x"2A",x"D4",x"40",x"EB",x"CD",x"C6",
x"29",x"CD",x"C6",x"29",x"21",x"49",x"23",x"E3",x"E5",x"C3",x"84",x"28",x"E1",x"E3",
x"7E",x"23",x"4E",x"23",x"46",x"6F",x"2C",x"2D",x"C8",x"0A",x"12",x"03",x"13",x"18",
x"F8",x"CD",x"F4",x"0A",x"2A",x"21",x"41",x"EB",x"CD",x"F5",x"29",x"EB",x"C0",x"D5",
x"50",x"59",x"1B",x"4E",x"2A",x"D6",x"40",x"DF",x"20",x"05",x"47",x"09",x"22",x"D6",
x"40",x"E1",x"C9",x"2A",x"B3",x"40",x"2B",x"46",x"2B",x"4E",x"2B",x"DF",x"C0",x"22",
x"B3",x"40",x"C9",x"01",x"F8",x"27",x"C5",x"CD",x"D7",x"29",x"AF",x"57",x"7E",x"B7",
x"C9",x"01",x"F8",x"27",x"C5",x"CD",x"07",x"2A",x"CA",x"4A",x"1E",x"23",x"5E",x"23",
x"56",x"1A",x"C9",x"3E",x"01",x"CD",x"57",x"28",x"CD",x"1F",x"2B",x"2A",x"D4",x"40",
x"73",x"C1",x"C3",x"84",x"28",x"D7",x"CF",x"28",x"CD",x"1C",x"2B",x"D5",x"CF",x"2C",
x"CD",x"37",x"23",x"CF",x"29",x"E3",x"E5",x"E7",x"28",x"05",x"CD",x"1F",x"2B",x"18",
x"03",x"CD",x"13",x"2A",x"D1",x"F5",x"F5",x"7B",x"CD",x"57",x"28",x"5F",x"F1",x"1C",
x"1D",x"28",x"D4",x"2A",x"D4",x"40",x"77",x"23",x"1D",x"20",x"FB",x"18",x"CA",x"CD",
x"DF",x"2A",x"AF",x"E3",x"4F",x"3E",x"E5",x"E5",x"7E",x"B8",x"38",x"02",x"78",x"11",
x"0E",x"00",x"C5",x"CD",x"BF",x"28",x"C1",x"E1",x"E5",x"23",x"46",x"23",x"66",x"68",
x"06",x"00",x"09",x"44",x"4D",x"CD",x"5A",x"28",x"6F",x"CD",x"CE",x"29",x"D1",x"CD",
x"DE",x"29",x"C3",x"84",x"28",x"CD",x"DF",x"2A",x"D1",x"D5",x"1A",x"90",x"18",x"CB",
x"EB",x"7E",x"CD",x"E2",x"2A",x"04",x"05",x"CA",x"4A",x"1E",x"C5",x"1E",x"FF",x"FE",
x"29",x"28",x"05",x"CF",x"2C",x"CD",x"1C",x"2B",x"CF",x"29",x"F1",x"E3",x"01",x"69",
x"2A",x"C5",x"3D",x"BE",x"06",x"00",x"D0",x"4F",x"7E",x"91",x"BB",x"47",x"D8",x"43",
x"C9",x"CD",x"07",x"2A",x"CA",x"F8",x"27",x"5F",x"23",x"7E",x"23",x"66",x"6F",x"E5",
x"19",x"46",x"72",x"E3",x"C5",x"7E",x"CD",x"65",x"0E",x"C1",x"E1",x"70",x"C9",x"EB",
x"CF",x"29",x"C1",x"D1",x"C5",x"43",x"C9",x"FE",x"7A",x"C2",x"97",x"19",x"C3",x"D9",
x"41",x"CD",x"1F",x"2B",x"32",x"94",x"40",x"CD",x"93",x"40",x"C3",x"F8",x"27",x"CD",
x"0E",x"2B",x"C3",x"96",x"40",x"D7",x"CD",x"37",x"23",x"E5",x"CD",x"7F",x"0A",x"EB",
x"E1",x"7A",x"B7",x"C9",x"CD",x"1C",x"2B",x"32",x"94",x"40",x"32",x"97",x"40",x"CF",
x"2C",x"18",x"01",x"D7",x"CD",x"37",x"23",x"CD",x"05",x"2B",x"C2",x"4A",x"1E",x"2B",
x"D7",x"7B",x"C9",x"3E",x"01",x"32",x"9C",x"40",x"C1",x"CD",x"10",x"1B",x"C5",x"21",
x"FF",x"FF",x"22",x"A2",x"40",x"E1",x"D1",x"4E",x"23",x"46",x"23",x"78",x"B1",x"CA",
x"19",x"1A",x"CD",x"DF",x"41",x"CD",x"9B",x"1D",x"C5",x"4E",x"23",x"46",x"23",x"C5",
x"E3",x"EB",x"DF",x"C1",x"DA",x"18",x"1A",x"E3",x"E5",x"C5",x"EB",x"22",x"EC",x"40",
x"CD",x"AF",x"0F",x"3E",x"20",x"E1",x"CD",x"2A",x"03",x"CD",x"7E",x"2B",x"2A",x"A7",
x"40",x"CD",x"75",x"2B",x"CD",x"FE",x"20",x"18",x"BE",x"7E",x"B7",x"C8",x"CD",x"2A",
x"03",x"23",x"18",x"F7",x"E5",x"2A",x"A7",x"40",x"44",x"4D",x"E1",x"16",x"FF",x"18",
x"03",x"03",x"15",x"C8",x"7E",x"B7",x"23",x"02",x"C8",x"F2",x"89",x"2B",x"FE",x"FB",
x"20",x"08",x"0B",x"0B",x"0B",x"0B",x"14",x"14",x"14",x"14",x"FE",x"95",x"CC",x"24",
x"0B",x"D6",x"7F",x"E5",x"5F",x"21",x"50",x"16",x"7E",x"B7",x"23",x"F2",x"AC",x"2B",
x"1D",x"20",x"F7",x"E6",x"7F",x"02",x"03",x"15",x"CA",x"D8",x"28",x"7E",x"23",x"B7",
x"F2",x"B7",x"2B",x"E1",x"18",x"C6",x"CD",x"10",x"1B",x"D1",x"C5",x"C5",x"CD",x"2C",
x"1B",x"30",x"05",x"54",x"5D",x"E3",x"E5",x"DF",x"D2",x"4A",x"1E",x"21",x"29",x"19",
x"CD",x"A7",x"28",x"C1",x"21",x"E8",x"1A",x"E3",x"EB",x"2A",x"F9",x"40",x"1A",x"02",
x"03",x"13",x"DF",x"20",x"F9",x"60",x"69",x"22",x"F9",x"40",x"C9",x"CD",x"84",x"02",
x"CD",x"37",x"23",x"E5",x"CD",x"13",x"2A",x"3E",x"D3",x"CD",x"64",x"02",x"CD",x"61",
x"02",x"1A",x"CD",x"64",x"02",x"2A",x"A4",x"40",x"EB",x"2A",x"F9",x"40",x"1A",x"13",
x"CD",x"64",x"02",x"DF",x"20",x"F8",x"CD",x"F8",x"01",x"E1",x"C9",x"CD",x"93",x"02",
x"7E",x"D6",x"B2",x"28",x"02",x"AF",x"01",x"2F",x"23",x"F5",x"2B",x"D7",x"3E",x"00",
x"28",x"07",x"CD",x"37",x"23",x"CD",x"13",x"2A",x"1A",x"6F",x"F1",x"B7",x"67",x"22",
x"21",x"41",x"CC",x"4D",x"1B",x"2A",x"21",x"41",x"EB",x"06",x"03",x"CD",x"35",x"02",
x"D6",x"D3",x"20",x"F7",x"10",x"F7",x"CD",x"35",x"02",x"1C",x"1D",x"28",x"03",x"BB",
x"20",x"37",x"2A",x"A4",x"40",x"06",x"03",x"CD",x"35",x"02",x"5F",x"96",x"A2",x"20",
x"21",x"73",x"CD",x"6C",x"19",x"7E",x"B7",x"23",x"20",x"ED",x"CD",x"2C",x"02",x"10",
x"EA",x"22",x"F9",x"40",x"21",x"29",x"19",x"CD",x"A7",x"28",x"CD",x"F8",x"01",x"2A",
x"A4",x"40",x"E5",x"C3",x"E8",x"1A",x"21",x"A5",x"2C",x"CD",x"A7",x"28",x"C3",x"18",
x"1A",x"32",x"3E",x"3C",x"06",x"03",x"CD",x"35",x"02",x"B7",x"20",x"F8",x"10",x"F8",
x"CD",x"96",x"02",x"18",x"A2",x"42",x"41",x"44",x"0D",x"00",x"CD",x"7F",x"0A",x"7E",
x"C3",x"F8",x"27",x"CD",x"02",x"2B",x"D5",x"CF",x"2C",x"CD",x"1C",x"2B",x"D1",x"12",
x"C9",x"CD",x"38",x"23",x"CD",x"F4",x"0A",x"CF",x"3B",x"EB",x"2A",x"21",x"41",x"18",
x"08",x"3A",x"DE",x"40",x"B7",x"28",x"0C",x"D1",x"EB",x"E5",x"AF",x"32",x"DE",x"40",
x"BA",x"F5",x"D5",x"46",x"B0",x"CA",x"4A",x"1E",x"23",x"4E",x"23",x"66",x"69",x"18",
x"1C",x"58",x"E5",x"0E",x"02",x"7E",x"23",x"FE",x"25",x"CA",x"17",x"2E",x"FE",x"20",
x"20",x"03",x"0C",x"10",x"F2",x"E1",x"43",x"3E",x"25",x"CD",x"49",x"2E",x"CD",x"2A",
x"03",x"AF",x"5F",x"57",x"CD",x"49",x"2E",x"57",x"7E",x"23",x"FE",x"21",x"CA",x"14",
x"2E",x"FE",x"23",x"28",x"37",x"05",x"CA",x"FE",x"2D",x"FE",x"2B",x"3E",x"08",x"28",
x"E7",x"2B",x"7E",x"23",x"FE",x"2E",x"28",x"40",x"FE",x"25",x"28",x"BD",x"BE",x"20",
x"D0",x"FE",x"24",x"28",x"14",x"FE",x"2A",x"20",x"C8",x"78",x"FE",x"02",x"23",x"38",
x"03",x"7E",x"FE",x"24",x"3E",x"20",x"20",x"07",x"05",x"1C",x"FE",x"AF",x"C6",x"10",
x"23",x"1C",x"82",x"57",x"1C",x"0E",x"00",x"05",x"28",x"47",x"7E",x"23",x"FE",x"2E",
x"28",x"18",x"FE",x"23",x"28",x"F0",x"FE",x"2C",x"20",x"1A",x"7A",x"F6",x"40",x"57",
x"18",x"E6",x"7E",x"FE",x"23",x"3E",x"2E",x"20",x"90",x"0E",x"01",x"23",x"0C",x"05",
x"28",x"25",x"7E",x"23",x"FE",x"23",x"28",x"F6",x"D5",x"11",x"97",x"2D",x"D5",x"54",
x"5D",x"FE",x"5B",x"C0",x"BE",x"C0",x"23",x"BE",x"C0",x"23",x"BE",x"C0",x"23",x"78",
x"D6",x"04",x"D8",x"D1",x"D1",x"47",x"14",x"23",x"CA",x"EB",x"D1",x"7A",x"2B",x"1C",
x"E6",x"08",x"20",x"15",x"1D",x"78",x"B7",x"28",x"10",x"7E",x"D6",x"2D",x"28",x"06",
x"FE",x"FE",x"20",x"07",x"3E",x"08",x"C6",x"04",x"82",x"57",x"05",x"E1",x"F1",x"28",
x"50",x"C5",x"D5",x"CD",x"37",x"23",x"D1",x"C1",x"C5",x"E5",x"43",x"78",x"81",x"FE",
x"19",x"D2",x"4A",x"1E",x"7A",x"F6",x"80",x"CD",x"BE",x"0F",x"CD",x"A7",x"28",x"E1",
x"2B",x"D7",x"37",x"28",x"0D",x"32",x"DE",x"40",x"FE",x"3B",x"28",x"05",x"FE",x"2C",
x"C2",x"97",x"19",x"D7",x"C1",x"EB",x"E1",x"E5",x"F5",x"D5",x"7E",x"90",x"23",x"4E",
x"23",x"66",x"69",x"16",x"00",x"5F",x"19",x"78",x"B7",x"C2",x"03",x"2D",x"18",x"06",
x"CD",x"49",x"2E",x"CD",x"2A",x"03",x"E1",x"F1",x"C2",x"CB",x"2C",x"DC",x"FE",x"20",
x"E3",x"CD",x"DD",x"29",x"E1",x"C3",x"69",x"21",x"0E",x"01",x"3E",x"F1",x"05",x"CD",
x"49",x"2E",x"E1",x"F1",x"28",x"E9",x"C5",x"CD",x"37",x"23",x"CD",x"F4",x"0A",x"C1",
x"C5",x"E5",x"2A",x"21",x"41",x"41",x"0E",x"00",x"C5",x"CD",x"68",x"2A",x"CD",x"AA",
x"28",x"2A",x"21",x"41",x"F1",x"96",x"47",x"3E",x"20",x"04",x"05",x"CA",x"D3",x"2D",
x"CD",x"2A",x"03",x"18",x"F7",x"F5",x"7A",x"B7",x"3E",x"2B",x"C4",x"2A",x"03",x"F1",
x"C9",x"32",x"9A",x"40",x"2A",x"EA",x"40",x"B4",x"A5",x"3C",x"EB",x"C8",x"18",x"04",
x"CD",x"4F",x"1E",x"C0",x"E1",x"EB",x"22",x"EC",x"40",x"EB",x"CD",x"2C",x"1B",x"D2",
x"D9",x"1E",x"60",x"69",x"23",x"23",x"4E",x"23",x"46",x"23",x"C5",x"CD",x"7E",x"2B",
x"E1",x"E5",x"CD",x"AF",x"0F",x"3E",x"20",x"CD",x"2A",x"03",x"2A",x"A7",x"40",x"3E",
x"0E",x"CD",x"2A",x"03",x"E5",x"0E",x"FF",x"0C",x"7E",x"B7",x"23",x"20",x"FA",x"E1",
x"47",x"16",x"00",x"CD",x"84",x"03",x"D6",x"30",x"38",x"0E",x"FE",x"0A",x"30",x"0A",
x"5F",x"7A",x"07",x"07",x"82",x"07",x"83",x"57",x"18",x"EB",x"E5",x"21",x"99",x"2E",
x"E3",x"15",x"14",x"C2",x"BB",x"2E",x"14",x"FE",x"D8",x"CA",x"D2",x"2F",x"FE",x"DD",
x"CA",x"E0",x"2F",x"FE",x"F0",x"28",x"41",x"FE",x"31",x"38",x"02",x"D6",x"20",x"FE",
x"21",x"CA",x"F6",x"2F",x"FE",x"1C",x"CA",x"40",x"2F",x"FE",x"23",x"28",x"3F",x"FE",
x"19",x"CA",x"7D",x"2F",x"FE",x"14",x"CA",x"4A",x"2F",x"FE",x"13",x"CA",x"65",x"2F",
x"FE",x"15",x"CA",x"E3",x"2F",x"FE",x"28",x"CA",x"78",x"2F",x"FE",x"1B",x"28",x"1C",
x"FE",x"18",x"CA",x"75",x"2F",x"FE",x"11",x"C0",x"C1",x"D1",x"CD",x"FE",x"20",x"C3",
x"65",x"2E",x"7E",x"B7",x"C8",x"04",x"CD",x"2A",x"03",x"23",x"15",x"20",x"F5",x"C9",
x"E5",x"21",x"5F",x"2F",x"E3",x"37",x"F5",x"CD",x"84",x"03",x"5F",x"F1",x"F5",x"DC",
x"5F",x"2F",x"7E",x"B7",x"CA",x"3E",x"2F",x"CD",x"2A",x"03",x"F1",x"F5",x"DC",x"A1",
x"2F",x"38",x"02",x"23",x"04",x"7E",x"BB",x"20",x"EB",x"15",x"20",x"E8",x"F1",x"C9",
x"CD",x"75",x"2B",x"CD",x"FE",x"20",x"C1",x"C3",x"7C",x"2E",x"7E",x"B7",x"C8",x"3E",
x"21",x"CD",x"2A",x"03",x"7E",x"B7",x"28",x"09",x"CD",x"2A",x"03",x"CD",x"A1",x"2F",
x"15",x"20",x"F3",x"3E",x"21",x"CD",x"2A",x"03",x"C9",x"7E",x"B7",x"C8",x"CD",x"84",
x"03",x"77",x"CD",x"2A",x"03",x"23",x"04",x"15",x"20",x"F1",x"C9",x"36",x"00",x"48",
x"16",x"FF",x"CD",x"0A",x"2F",x"CD",x"84",x"03",x"B7",x"CA",x"7D",x"2F",x"FE",x"08",
x"28",x"0A",x"FE",x"0D",x"CA",x"E0",x"2F",x"FE",x"1B",x"C8",x"20",x"1E",x"3E",x"08",
x"05",x"04",x"28",x"1F",x"CD",x"2A",x"03",x"2B",x"05",x"11",x"7D",x"2F",x"D5",x"E5",
x"0D",x"7E",x"B7",x"37",x"CA",x"90",x"08",x"23",x"7E",x"2B",x"77",x"23",x"18",x"F3",
x"F5",x"79",x"FE",x"FF",x"38",x"03",x"F1",x"18",x"C4",x"90",x"0C",x"04",x"C5",x"EB",
x"6F",x"26",x"00",x"19",x"44",x"4D",x"23",x"CD",x"58",x"19",x"C1",x"F1",x"77",x"CD",
x"2A",x"03",x"23",x"C3",x"7D",x"2F",x"78",x"B7",x"C8",x"05",x"2B",x"3E",x"08",x"CD",
x"2A",x"03",x"15",x"20",x"F3",x"C9",x"CD",x"75",x"2B",x"CD",x"FE",x"20",x"C1",x"D1",
x"7A",x"A3",x"3C",x"2A",x"A7",x"40",x"2B",x"C8",x"37",x"23",x"F5",x"C3",x"98",x"1A",
x"C1",x"D1",x"C3",x"19",x"1A",x"DE",x"C3",x"C3",x"44",x"B2",
x"CD",x"5C",x"30",x"C3",x"21",x"30",x"21",x"47",x"31",x"18",x"07",x"CD",x"5C",x"30",
x"3E",x"10",x"18",x"10",x"22",x"1E",x"40",x"21",x"D4",x"33",x"22",x"04",x"40",x"CD",
x"61",x"1B",x"C3",x"19",x"1A",x"AF",x"FD",x"77",x"06",x"FD",x"E5",x"E1",x"06",x"05",
x"AF",x"23",x"77",x"10",x"FC",x"21",x"40",x"30",x"CD",x"C9",x"01",x"CD",x"A7",x"28",
x"21",x"78",x"30",x"22",x"16",x"40",x"18",x"C6",x"4E",x"45",x"57",x"20",x"4B",x"45",
x"59",x"42",x"4F",x"41",x"52",x"44",x"20",x"52",x"4F",x"55",x"54",x"49",x"4E",x"45",
x"20",x"45",x"4E",x"41",x"42",x"4C",x"45",x"00",x"2A",x"B1",x"40",x"11",x"FA",x"FF",
x"19",x"22",x"B1",x"40",x"22",x"49",x"40",x"22",x"1B",x"40",x"11",x"CE",x"FF",x"19",
x"22",x"A0",x"40",x"FD",x"2A",x"1B",x"40",x"C9",x"FD",x"E5",x"CD",x"80",x"30",x"FD",
x"E1",x"C9",x"FD",x"2A",x"1B",x"40",x"21",x"36",x"40",x"01",x"80",x"38",x"0A",x"E6",
x"01",x"28",x"14",x"0E",x"40",x"0A",x"E6",x"04",x"28",x"0D",x"0A",x"E6",x"04",x"20",
x"FB",x"FD",x"7E",x"06",x"EE",x"10",x"FD",x"77",x"06",x"FD",x"7E",x"05",x"A7",x"28",
x"08",x"5F",x"FD",x"4E",x"03",x"0A",x"A3",x"20",x"47",x"3A",x"22",x"40",x"A7",x"28",
x"13",x"FD",x"7E",x"06",x"A7",x"20",x"0D",x"FD",x"34",x"02",x"20",x"08",x"ED",x"5B",
x"20",x"40",x"1A",x"EE",x"D0",x"12",x"AF",x"FD",x"77",x"05",x"0E",x"01",x"16",x"00",
x"0A",x"5F",x"AE",x"73",x"A3",x"20",x"08",x"14",x"2C",x"CB",x"01",x"F2",x"D2",x"30",
x"C9",x"5F",x"C5",x"01",x"00",x"06",x"CD",x"60",x"00",x"C1",x"0A",x"A3",x"C8",x"FD",
x"77",x"05",x"FD",x"71",x"03",x"FD",x"70",x"04",x"18",x"6D",x"FD",x"7E",x"04",x"A7",
x"20",x"0E",x"C5",x"01",x"00",x"0A",x"CD",x"60",x"00",x"C1",x"0A",x"A3",x"28",x"C0",
x"18",x"28",x"21",x"00",x"4C",x"E5",x"C5",x"21",x"36",x"40",x"0E",x"01",x"0A",x"5F",
x"AE",x"A3",x"20",x"23",x"2C",x"CB",x"01",x"F2",x"16",x"31",x"C1",x"FD",x"5E",x"05",
x"0A",x"A3",x"28",x"16",x"E1",x"2B",x"CB",x"74",x"20",x"DF",x"AF",x"FD",x"77",x"04",
x"16",x"00",x"CB",x"41",x"20",x"2B",x"CB",x"19",x"14",x"18",x"F7",x"C1",x"E1",x"21",
x"36",x"40",x"C3",x"CA",x"30",x"DD",x"6E",x"03",x"DD",x"66",x"04",x"DA",x"9A",x"04",
x"DD",x"7E",x"05",x"B7",x"28",x"01",x"77",x"79",x"FE",x"20",x"DA",x"06",x"05",x"FE",
x"80",x"D2",x"A6",x"04",x"C3",x"7D",x"04",x"E5",x"21",x"6D",x"31",x"E3",x"C3",x"FB",
x"03",x"FE",x"10",x"28",x"01",x"C9",x"DB",x"FD",x"E6",x"F0",x"FE",x"30",x"20",x"2A",
x"21",x"00",x"3C",x"7D",x"E6",x"3F",x"3E",x"0D",x"CC",x"3B",x"00",x"7E",x"CB",x"7F",
x"28",x"02",x"E6",x"BF",x"CB",x"74",x"23",x"20",x"05",x"CD",x"3B",x"00",x"18",x"E7",
x"06",x"06",x"3E",x"20",x"CD",x"3B",x"00",x"3E",x"0D",x"CD",x"3B",x"00",x"10",x"F4",
x"AF",x"C9",x"E3",x"22",x"FE",x"41",x"E3",x"ED",x"73",x"FC",x"41",x"31",x"FC",x"41",
x"08",x"D9",x"E5",x"D5",x"C5",x"F5",x"08",x"D9",x"E5",x"D5",x"C5",x"F5",x"DD",x"E5",
x"FD",x"E5",x"ED",x"7B",x"FC",x"41",x"CD",x"C9",x"01",x"CD",x"34",x"32",x"CD",x"49",
x"00",x"CD",x"3A",x"03",x"FE",x"44",x"28",x"19",x"FE",x"4D",x"28",x"4D",x"FE",x"52",
x"28",x"4E",x"FE",x"42",x"20",x"06",x"CD",x"61",x"1B",x"C3",x"19",x"1A",x"FE",x"47",
x"CC",x"EB",x"32",x"18",x"D7",x"CD",x"92",x"33",x"FE",x"58",x"28",x"D0",x"CD",x"C9",
x"01",x"CD",x"69",x"32",x"3E",x"3E",x"CD",x"3A",x"03",x"06",x"10",x"7E",x"CD",x"73",
x"33",x"3E",x"20",x"CD",x"3A",x"03",x"23",x"10",x"F4",x"3E",x"0D",x"CD",x"3A",x"03",
x"CD",x"49",x"00",x"FE",x"0A",x"28",x"DE",x"FE",x"5B",x"20",x"A7",x"11",x"20",x"00",
x"B7",x"ED",x"52",x"18",x"D2",x"CD",x"72",x"32",x"18",x"9A",x"CD",x"C9",x"01",x"CD",
x"BD",x"32",x"18",x"92",x"FD",x"21",x"E8",x"41",x"21",x"98",x"32",x"06",x"0C",x"C5",
x"CD",x"4E",x"32",x"3E",x"0D",x"CD",x"3A",x"03",x"C1",x"FD",x"23",x"FD",x"23",x"10",
x"F0",x"C9",x"06",x"03",x"7E",x"CD",x"3A",x"03",x"23",x"10",x"F9",x"3E",x"3D",x"CD",
x"3A",x"03",x"FD",x"7E",x"01",x"CD",x"73",x"33",x"FD",x"7E",x"00",x"CD",x"73",x"33",
x"C9",x"7C",x"CD",x"73",x"33",x"7D",x"CD",x"73",x"33",x"C9",x"CD",x"92",x"33",x"FE",
x"58",x"C8",x"CD",x"C9",x"01",x"CD",x"69",x"32",x"3E",x"3E",x"CD",x"3A",x"03",x"7E",
x"CD",x"73",x"33",x"3E",x"2D",x"CD",x"3A",x"03",x"CD",x"9B",x"33",x"70",x"3E",x"0D",
x"CD",x"3A",x"03",x"23",x"18",x"E3",x"49",x"59",x"20",x"49",x"58",x"20",x"41",x"46",
x"20",x"42",x"43",x"20",x"44",x"45",x"20",x"48",x"4C",x"20",x"41",x"46",x"27",x"42",
x"43",x"27",x"44",x"45",x"27",x"48",x"4C",x"27",x"53",x"50",x"20",x"50",x"43",x"20",
x"00",x"21",x"98",x"32",x"FD",x"21",x"E8",x"41",x"06",x"0C",x"C5",x"CD",x"4E",x"32",
x"3E",x"2F",x"CD",x"3A",x"03",x"E5",x"CD",x"92",x"33",x"FE",x"58",x"28",x"06",x"FD",
x"75",x"00",x"FD",x"74",x"01",x"FD",x"23",x"FD",x"23",x"E1",x"3E",x"0D",x"CD",x"3A",
x"03",x"C1",x"10",x"DC",x"C9",x"CD",x"9B",x"33",x"60",x"CD",x"9B",x"33",x"68",x"22",
x"FE",x"41",x"CD",x"49",x"00",x"FE",x"2C",x"28",x"09",x"FE",x"0D",x"28",x"22",x"FE",
x"58",x"C8",x"18",x"F0",x"CD",x"3A",x"03",x"CD",x"92",x"33",x"FE",x"58",x"C8",x"E5",
x"11",x"00",x"42",x"01",x"03",x"00",x"ED",x"B0",x"E1",x"11",x"47",x"33",x"3E",x"CD",
x"77",x"23",x"73",x"23",x"72",x"ED",x"7B",x"FC",x"41",x"2A",x"FE",x"41",x"E5",x"ED",
x"73",x"FC",x"41",x"31",x"E8",x"41",x"FD",x"E1",x"DD",x"E1",x"F1",x"C1",x"D1",x"E1",
x"08",x"D9",x"F1",x"C1",x"D1",x"E1",x"08",x"D9",x"ED",x"7B",x"FC",x"41",x"C9",x"E3",
x"2B",x"2B",x"2B",x"22",x"FE",x"41",x"32",x"03",x"42",x"ED",x"53",x"04",x"42",x"78",
x"32",x"06",x"42",x"11",x"00",x"42",x"EB",x"01",x"03",x"00",x"ED",x"B0",x"EB",x"ED",
x"5B",x"04",x"42",x"3A",x"06",x"42",x"47",x"3A",x"03",x"42",x"21",x"AB",x"31",x"E3",
x"C9",x"4F",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"CD",x"86",x"33",x"79",
x"E6",x"0F",x"CD",x"86",x"33",x"C9",x"C6",x"30",x"FE",x"3A",x"38",x"02",x"C6",x"07",
x"CD",x"3A",x"03",x"C9",x"CD",x"9B",x"33",x"60",x"CD",x"9B",x"33",x"68",x"C9",x"CD",
x"B5",x"33",x"CB",x"27",x"CB",x"27",x"CB",x"27",x"CB",x"27",x"47",x"79",x"CD",x"3A",
x"03",x"CD",x"B5",x"33",x"80",x"47",x"79",x"CD",x"3A",x"03",x"C9",x"CD",x"49",x"00",
x"FE",x"58",x"20",x"05",x"E3",x"E1",x"E3",x"E1",x"C9",x"4F",x"D6",x"30",x"38",x"EF",
x"FE",x"0A",x"D8",x"D6",x"11",x"38",x"E8",x"C6",x"0A",x"FE",x"10",x"D8",x"18",x"E1",
x"E3",x"3E",x"1D",x"BC",x"20",x"03",x"3E",x"5B",x"BD",x"E3",x"C2",x"78",x"1D",x"CD",
x"78",x"1D",x"F5",x"E5",x"FE",x"52",x"20",x"07",x"23",x"7E",x"FE",x"45",x"CA",x"6D",
x"34",x"E1",x"F1",x"C9",x"D5",x"22",x"21",x"41",x"01",x"00",x"00",x"2A",x"A7",x"40",
x"E5",x"CD",x"2F",x"13",x"E1",x"06",x"05",x"7E",x"D6",x"30",x"20",x"05",x"23",x"10",
x"F8",x"2B",x"04",x"D1",x"C9",x"FD",x"23",x"FD",x"23",x"FD",x"23",x"FD",x"23",x"C9",
x"23",x"7E",x"B7",x"C8",x"FE",x"8D",x"28",x"0C",x"FE",x"91",x"28",x"08",x"FE",x"CA",
x"28",x"04",x"FE",x"95",x"20",x"EC",x"A7",x"C9",x"ED",x"5B",x"A7",x"40",x"D5",x"06",
x"00",x"7E",x"FE",x"20",x"28",x"0B",x"FE",x"30",x"38",x"0A",x"FE",x"3A",x"30",x"06",
x"04",x"12",x"13",x"23",x"18",x"ED",x"AF",x"12",x"D1",x"04",x"05",x"C9",x"C5",x"78",
x"99",x"28",x"10",x"05",x"28",x"08",x"0D",x"20",x"F6",x"CD",x"CD",x"35",x"18",x"05",
x"41",x"05",x"CD",x"AC",x"35",x"C1",x"1A",x"77",x"13",x"23",x"10",x"FA",x"C9",x"23",
x"11",x"0A",x"00",x"ED",x"53",x"E2",x"40",x"ED",x"53",x"E4",x"40",x"7E",x"A7",x"28",
x"22",x"FE",x"2C",x"28",x"11",x"CD",x"5A",x"1E",x"4F",x"7A",x"B3",x"28",x"13",x"79",
x"ED",x"53",x"E2",x"40",x"FE",x"2C",x"20",x"0D",x"23",x"CD",x"5A",x"1E",x"ED",x"53",
x"E4",x"40",x"7A",x"B3",x"CA",x"97",x"19",x"FD",x"2A",x"F9",x"40",x"11",x"00",x"01",
x"FD",x"19",x"FD",x"E5",x"2A",x"A4",x"40",x"E5",x"7E",x"23",x"B6",x"CA",x"FE",x"34",
x"23",x"23",x"CD",x"1A",x"34",x"23",x"28",x"F2",x"CD",x"30",x"34",x"2B",x"28",x"F4",
x"23",x"E5",x"D5",x"FD",x"E5",x"D1",x"2A",x"B1",x"40",x"ED",x"52",x"DA",x"7A",x"19",
x"11",x"04",x"00",x"ED",x"52",x"DA",x"7A",x"19",x"FD",x"70",x"00",x"E1",x"CD",x"5A",
x"1E",x"FD",x"73",x"01",x"FD",x"72",x"02",x"FD",x"36",x"03",x"00",x"CD",x"11",x"34",
x"E1",x"2B",x"23",x"7E",x"FE",x"20",x"28",x"FA",x"FE",x"2C",x"28",x"03",x"2B",x"18",
x"BB",x"23",x"18",x"BE",x"FD",x"36",x"00",x"FF",x"E1",x"FD",x"E1",x"ED",x"5B",x"E2",
x"40",x"D5",x"FD",x"E5",x"E5",x"D5",x"CD",x"C2",x"09",x"7A",x"B3",x"28",x"41",x"EB",
x"D1",x"FD",x"E5",x"FD",x"7E",x"00",x"3C",x"28",x"21",x"FD",x"7E",x"03",x"B7",x"20",
x"16",x"FD",x"7E",x"01",x"B9",x"20",x"10",x"FD",x"7E",x"02",x"B8",x"20",x"0A",x"FD",
x"73",x"01",x"FD",x"72",x"02",x"FD",x"36",x"03",x"01",x"CD",x"11",x"34",x"18",x"D9",
x"FD",x"E1",x"E5",x"2A",x"E4",x"40",x"19",x"DA",x"7A",x"19",x"EB",x"21",x"F8",x"FF",
x"ED",x"52",x"DA",x"7A",x"19",x"E1",x"18",x"B7",x"D1",x"E1",x"FD",x"E1",x"D1",x"7E",
x"23",x"B6",x"CA",x"83",x"2C",x"23",x"73",x"23",x"72",x"CD",x"1A",x"34",x"23",x"20",
x"09",x"E5",x"2A",x"E4",x"40",x"19",x"EB",x"E1",x"18",x"E7",x"E5",x"D5",x"CD",x"30",
x"34",x"D1",x"E1",x"2B",x"28",x"E7",x"23",x"7E",x"FE",x"20",x"28",x"FA",x"D5",x"E5",
x"FD",x"6E",x"01",x"FD",x"66",x"02",x"CD",x"F4",x"33",x"FD",x"4E",x"00",x"CD",x"11",
x"34",x"EB",x"E1",x"CD",x"50",x"34",x"D1",x"2B",x"23",x"7E",x"FE",x"20",x"28",x"FA",
x"FE",x"2C",x"28",x"03",x"2B",x"18",x"BC",x"23",x"18",x"C8",x"D5",x"C5",x"E5",x"E5",
x"D1",x"D5",x"D5",x"2A",x"F9",x"40",x"E5",x"2B",x"13",x"10",x"FC",x"22",x"F9",x"40",
x"E1",x"C1",x"ED",x"42",x"23",x"E5",x"C1",x"E1",x"EB",x"ED",x"B0",x"E1",x"C1",x"D1",
x"C9",x"D5",x"C5",x"E5",x"2A",x"F9",x"40",x"E5",x"D1",x"23",x"10",x"FD",x"22",x"F9",
x"40",x"C1",x"C5",x"E5",x"B7",x"ED",x"42",x"E5",x"C1",x"03",x"E1",x"EB",x"ED",x"B8",
x"E1",x"C1",x"D1",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",

others => x"ff"
  );

signal  do : std_logic_vector(7 downto 0);

begin

  process(CLK)
  begin
    if rising_edge(CLK) then
	   do <= myROM(conv_integer(A));
	 end if;
  end process;  
  DOUT <= do;
  
end Behavioral;
