-------------------------------------------------------------------------------
--
-- The BUS unit.
-- Implements the BUS port logic.
--
-- $Id: db_bus-c.vhd,v 1.2 2005/06/11 10:08:43 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_db_bus_rtl_c0 of t48_db_bus is

  for rtl
  end for;

end t48_db_bus_rtl_c0;
