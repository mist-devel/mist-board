`timescale  1 ps / 1 ps
