module dongle (
	// cpu register interface
	input 		 clk,
	input 		 sel,
	input 		 cpu_as, // cpu_cycle && as
	input 		 uds,
	input 		 rw,
	input [14:0] 	 addr,
	output reg [7:0] dout,
		
	output 		 present
);

assign present = 1'b0;  // 0 = deactivate dongle

// ------------------------------------------------------------------------------------
// ------------------------------------ CUBASE 2 DONGLE -------------------------------
// ------------------------------------------------------------------------------------
reg [15:8] d;
reg [15:8] next_d;

// read
always @(sel, uds, rw, d) begin
	dout = 8'd0;
	if(sel && ~uds && rw)
		dout = d;
end

wire [8:1] a = addr[7:0];

// special addresses: 
// a[8:1] = 8'b11011000,0 -> 0x1b0     clear all
// a[8:1] = 8'bxxx00xx0,0 ->  a5+a4+a1 = 0 sets all, incl. $0c
   
// update register in the middle of the transfer
always @(negedge clk) begin
	if(cpu_as && ~uds) begin
      next_d[15] <= !(( a[8] & a[7] & !a[6] & a[5] & a[4] & !a[3] & !a[2] & !a[1]) | 
                 (!d[15] & !d[14] & !d[13] & !d[12] & !d[11] &  d[10] & !d[9]         & a[4]       ) | 
                 (          d[14]          &  d[12]          &  d[10]                        & a[1]) | 
                 (                   d[13] &                   !d[10]                 & a[4]       ) | 
                 (         !d[14]                            & !d[10]                        & a[1]) | 
                 ( d[15]                                     & !d[10]                 & a[4]       ) | 
                 (                           !d[12]          & !d[10]                        & a[1]) | 
                 (!d[8] & a[5] ));
      
      next_d[14] <= !(( a[8] & a[7] & !a[6] & a[5] & a[4] & !a[3] & !a[2] & !a[1]) | 
                 (!d[15] & !d[14] & !d[13] & !d[12] & !d[11] & !d[10] & !d[9] &  d[8] & a[4]       ) | 
                 (          d[14]          &  d[12]          &  d[10]         &  d[8]        & a[1]) | 
                 (                                             !d[10]         & !d[8]        & a[1]) | 
                 (                           !d[12]                           & !d[8]        & a[1]) | 
                 ( d[15]                                                      & !d[8] & a[4]       ) | 
                 (         !d[14]                                             & !d[8]        & a[1]) | 
                 (!d[15] & a[5] ));
      
      next_d[13] <= !(( a[8] & a[7] & !a[6] & a[5] & a[4] & !a[3] & !a[2] & !a[1]) | 
                 (d[15]&d[14]&d[13]&d[12]&d[11]&d[10]&d[8]&a[1]) | 
                 (!d[15]&!d[13]&d[11]&a[4]) | 
                 (d[13]&!d[11]&a[4]) | 
                 (!d[12]&!d[11]&a[1]) | 
                 (d[15]&!d[11]&a[4]) | 
                 (!d[14]&!d[11]&a[1]) | 
                 (!d[9]&a[5]));

      next_d[12] <= !(( a[8] & a[7] & !a[6] & a[5] & a[4] & !a[3] & !a[2] & !a[1]) |
                 (d[15]&d[14]&d[13]&d[12]&d[10]&d[8]&a[1]) | 
                 (!d[13]&!d[10]&a[1]) | 
                 (!d[15]&d[13]&a[4]) | 
                 (!d[13]&!d[12]&a[1]) | 
                 (d[15]&!d[13]&a[4]) |
                 (!d[14]&!d[13]&a[1]) |
                 (!d[11]&a[5]));
					  
     next_d[11] <= !(( a[8] & a[7] & !a[6] & a[5] & a[4] & !a[3] & !a[2] & !a[1]) |
                 (d[15]&d[14]&d[12]&d[10]&d[8]&a[1]) |
                 (!d[15]&!d[8]&a[1]) |
                 (!d[15]&!d[10]&a[1]) |
                 (!d[15]&!d[12]&a[1]) |
                 (!d[15]&!d[14]&a[1]) |
                 (d[15]&a[4]) |
                 (!d[13]&a[5]));

      next_d[10] <= !(( a[8] & a[7] & !a[6] & a[5] & a[4] & !a[3] & !a[2] & !a[1]) |
                 (d[15]&d[14]&d[13]&d[12]&d[11]&d[10]&d[9]&d[8]&a[1]) |
                 (!d[15]&!d[13]&!d[11]&d[9]&a[4]) |
                 (d[11]&!d[9]&a[4]) |
                 (d[13]&!d[9]&a[4]) |
                 (d[15]&!d[9]&a[4]) |
                 (!d[14]&!d[9]&a[1]) |
                 (!d[14]&a[5]));

      next_d[9] <= !(( a[8] & a[7] & !a[6] & a[5] & a[4] & !a[3] & !a[2] & !a[1]) |
                (!d[15]&d[14]&!d[13]&!d[11]&!d[9]&a[4]) |
                (!d[14]&d[9]&a[4]) |
                (!d[14]&d[11]&a[4]) |
                (!d[14]&d[13]&a[4]) |
                (d[15]&!d[14]&a[4]) |
                (d[14]&a[1]) |
                (!d[12]&a[5]));

      next_d[8] <= !(( a[8] & a[7] & !a[6] & a[5] & a[4] & !a[3] & !a[2] & !a[1]) |
                (!d[15]&!d[14]&!d[13]&d[12]&!d[11]&!d[9]&a[4]) |
                (d[14]&d[12]&a[1]) |
                (!d[12]&d[11]&a[4]) |
                (d[13]&!d[12]&a[4]) |
                (d[15]&!d[12]&a[4]) |
                (!d[14]&!d[12]&a[1]) |
                (!d[10]&a[5]));
					  
					  
	end
end

always @(posedge clk)
	d <= next_d;

endmodule