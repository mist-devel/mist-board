-------------------------------------------------------------------------------
--
-- $Id: clock_ctrl-c.vhd,v 1.2 2005/06/11 10:08:43 arniml Exp $
--
-- The clock control unit.
--
-------------------------------------------------------------------------------

configuration t48_clock_ctrl_rtl_c0 of t48_clock_ctrl is

  for rtl
  end for;

end t48_clock_ctrl_rtl_c0;
