-------------------------------------------------------------------------------
--
-- T8x48 ROM
--
-- $Id: t48_rom-struct-a.vhd,v 1.1.1.3 2006/11/26 10:07:52 arnim Exp $
--
-- Copyright (c) 2006 Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-- Redistribution and use in source and synthezised forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- Please report bugs to the author, but before you do so, please
-- make sure that this is not a derivative work and that
-- you have the latest version of this file.
--
-- The latest version of this file can be found at:
--      http://www.opencores.org/cvsweb.shtml/t48/
--
-------------------------------------------------------------------------------

architecture struct of t48_rom is

  component rom_t48
    port(
      Clk : in  std_logic;
      A   : in  std_logic_vector(9 downto 0);
      D   : out std_logic_vector(7 downto 0)
    );
  end component;

begin

  rom_b : rom_t48
    port map (
      Clk => clk_i,
      A   => rom_addr_i,
      D   => rom_data_o
    );

end struct;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t48_rom-struct-a.vhd,v $
-- Revision 1.1.1.3  2006/11/26 10:07:52  arnim
-- incremental import for release 1.0
--
-- Revision 1.3  2006/11/26 12:53:28  arniml
-- fix entity port names
--
-- Revision 1.2  2006/11/26 11:58:28  arniml
-- fix component name
--
-- Revision 1.1  2006/06/21 00:59:15  arniml
-- initial check-in
--
-------------------------------------------------------------------------------
