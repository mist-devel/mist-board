-------------------------------------------------------------------------------
--
-- The Port 2 unit.
-- Implements the Port 2 logic.
--
-- $Id: p2-c.vhd,v 1.2 2005/06/11 10:08:43 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_p2_rtl_c0 of t48_p2 is

  for rtl
  end for;

end t48_p2_rtl_c0;
