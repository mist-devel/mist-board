-------------------------------------------------------------------------------
--
-- The Port 1 unit.
-- Implements the Port 1 logic.
--
-- $Id: p1-c.vhd,v 1.2 2005/06/11 10:08:43 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_p1_rtl_c0 of t48_p1 is

  for rtl
  end for;

end t48_p1_rtl_c0;
