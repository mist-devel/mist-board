-------------------------------------------------------------------------------
--
-- Synthesizable model of TI's SN76489AN.
--
-- $Id: sn76489_clock_div-c.vhd,v 1.2 2005/10/10 22:12:38 arnim Exp $
--
-------------------------------------------------------------------------------

configuration sn76489_clock_div_rtl_c0 of sn76489_clock_div is

  for rtl
  end for;

end sn76489_clock_div_rtl_c0;
